magic
tech sky130A
magscale 1 2
timestamp 1764771510
<< viali >>
rect 6009 8041 6043 8075
rect 1409 7837 1443 7871
rect 3893 7837 3927 7871
rect 6101 7769 6135 7803
rect 1593 7701 1627 7735
rect 3985 7701 4019 7735
rect 6653 6817 6687 6851
rect 6101 6613 6135 6647
rect 5917 6273 5951 6307
rect 6193 6273 6227 6307
rect 5273 6205 5307 6239
rect 6009 6069 6043 6103
rect 5076 5865 5110 5899
rect 6561 5865 6595 5899
rect 1961 5729 1995 5763
rect 2053 5729 2087 5763
rect 4813 5729 4847 5763
rect 2145 5593 2179 5627
rect 2513 5525 2547 5559
rect 5089 5321 5123 5355
rect 6009 5321 6043 5355
rect 1777 5253 1811 5287
rect 5457 5185 5491 5219
rect 5549 5185 5583 5219
rect 6101 5185 6135 5219
rect 2053 5117 2087 5151
rect 2329 5117 2363 5151
rect 3801 5117 3835 5151
rect 4905 5117 4939 5151
rect 5641 5117 5675 5151
rect 1501 4981 1535 5015
rect 4353 4981 4387 5015
rect 1961 4777 1995 4811
rect 2789 4709 2823 4743
rect 3433 4641 3467 4675
rect 6101 4641 6135 4675
rect 6193 4641 6227 4675
rect 1777 4573 1811 4607
rect 2237 4573 2271 4607
rect 3249 4573 3283 4607
rect 3801 4505 3835 4539
rect 2053 4437 2087 4471
rect 3157 4437 3191 4471
rect 5089 4437 5123 4471
rect 5641 4437 5675 4471
rect 6009 4437 6043 4471
rect 2789 4233 2823 4267
rect 3893 4233 3927 4267
rect 5825 4165 5859 4199
rect 3341 4097 3375 4131
rect 3985 4097 4019 4131
rect 6101 4029 6135 4063
rect 3433 3689 3467 3723
rect 1685 3553 1719 3587
rect 4813 3485 4847 3519
rect 5273 3485 5307 3519
rect 1961 3417 1995 3451
rect 4629 3349 4663 3383
rect 5365 3349 5399 3383
rect 1869 3145 1903 3179
rect 3341 3145 3375 3179
rect 5733 3145 5767 3179
rect 3157 3077 3191 3111
rect 4445 3077 4479 3111
rect 3433 3009 3467 3043
rect 4077 3009 4111 3043
rect 3985 2805 4019 2839
rect 6009 2601 6043 2635
rect 6469 2533 6503 2567
rect 4261 2465 4295 2499
rect 4537 2329 4571 2363
rect 6653 2329 6687 2363
<< metal1 >>
rect 1104 8186 7084 8208
rect 1104 8134 1697 8186
rect 1749 8134 1761 8186
rect 1813 8134 1825 8186
rect 1877 8134 1889 8186
rect 1941 8134 1953 8186
rect 2005 8134 3192 8186
rect 3244 8134 3256 8186
rect 3308 8134 3320 8186
rect 3372 8134 3384 8186
rect 3436 8134 3448 8186
rect 3500 8134 4687 8186
rect 4739 8134 4751 8186
rect 4803 8134 4815 8186
rect 4867 8134 4879 8186
rect 4931 8134 4943 8186
rect 4995 8134 6182 8186
rect 6234 8134 6246 8186
rect 6298 8134 6310 8186
rect 6362 8134 6374 8186
rect 6426 8134 6438 8186
rect 6490 8134 7084 8186
rect 1104 8112 7084 8134
rect 5997 8075 6055 8081
rect 5997 8041 6009 8075
rect 6043 8072 6055 8075
rect 7742 8072 7748 8084
rect 6043 8044 7748 8072
rect 6043 8041 6055 8044
rect 5997 8035 6055 8041
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 3660 7840 3893 7868
rect 3660 7828 3666 7840
rect 3881 7837 3893 7840
rect 3927 7837 3939 7871
rect 3881 7831 3939 7837
rect 6086 7760 6092 7812
rect 6144 7760 6150 7812
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 2038 7732 2044 7744
rect 1627 7704 2044 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 3050 7692 3056 7744
rect 3108 7732 3114 7744
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3108 7704 3985 7732
rect 3108 7692 3114 7704
rect 3973 7701 3985 7704
rect 4019 7701 4031 7735
rect 3973 7695 4031 7701
rect 1104 7642 7156 7664
rect 1104 7590 2357 7642
rect 2409 7590 2421 7642
rect 2473 7590 2485 7642
rect 2537 7590 2549 7642
rect 2601 7590 2613 7642
rect 2665 7590 3852 7642
rect 3904 7590 3916 7642
rect 3968 7590 3980 7642
rect 4032 7590 4044 7642
rect 4096 7590 4108 7642
rect 4160 7590 5347 7642
rect 5399 7590 5411 7642
rect 5463 7590 5475 7642
rect 5527 7590 5539 7642
rect 5591 7590 5603 7642
rect 5655 7590 6842 7642
rect 6894 7590 6906 7642
rect 6958 7590 6970 7642
rect 7022 7590 7034 7642
rect 7086 7590 7098 7642
rect 7150 7590 7156 7642
rect 1104 7568 7156 7590
rect 1104 7098 7084 7120
rect 1104 7046 1697 7098
rect 1749 7046 1761 7098
rect 1813 7046 1825 7098
rect 1877 7046 1889 7098
rect 1941 7046 1953 7098
rect 2005 7046 3192 7098
rect 3244 7046 3256 7098
rect 3308 7046 3320 7098
rect 3372 7046 3384 7098
rect 3436 7046 3448 7098
rect 3500 7046 4687 7098
rect 4739 7046 4751 7098
rect 4803 7046 4815 7098
rect 4867 7046 4879 7098
rect 4931 7046 4943 7098
rect 4995 7046 6182 7098
rect 6234 7046 6246 7098
rect 6298 7046 6310 7098
rect 6362 7046 6374 7098
rect 6426 7046 6438 7098
rect 6490 7046 7084 7098
rect 1104 7024 7084 7046
rect 6086 6808 6092 6860
rect 6144 6848 6150 6860
rect 6546 6848 6552 6860
rect 6144 6820 6552 6848
rect 6144 6808 6150 6820
rect 6546 6808 6552 6820
rect 6604 6848 6610 6860
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 6604 6820 6653 6848
rect 6604 6808 6610 6820
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 5132 6616 6101 6644
rect 5132 6604 5138 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 6089 6607 6147 6613
rect 1104 6554 7156 6576
rect 1104 6502 2357 6554
rect 2409 6502 2421 6554
rect 2473 6502 2485 6554
rect 2537 6502 2549 6554
rect 2601 6502 2613 6554
rect 2665 6502 3852 6554
rect 3904 6502 3916 6554
rect 3968 6502 3980 6554
rect 4032 6502 4044 6554
rect 4096 6502 4108 6554
rect 4160 6502 5347 6554
rect 5399 6502 5411 6554
rect 5463 6502 5475 6554
rect 5527 6502 5539 6554
rect 5591 6502 5603 6554
rect 5655 6502 6842 6554
rect 6894 6502 6906 6554
rect 6958 6502 6970 6554
rect 7022 6502 7034 6554
rect 7086 6502 7098 6554
rect 7150 6502 7156 6554
rect 1104 6480 7156 6502
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6304 5963 6307
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 5951 6276 6193 6304
rect 5951 6273 5963 6276
rect 5905 6267 5963 6273
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 5258 6196 5264 6248
rect 5316 6196 5322 6248
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 5592 6072 6009 6100
rect 5592 6060 5598 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 5997 6063 6055 6069
rect 1104 6010 7084 6032
rect 1104 5958 1697 6010
rect 1749 5958 1761 6010
rect 1813 5958 1825 6010
rect 1877 5958 1889 6010
rect 1941 5958 1953 6010
rect 2005 5958 3192 6010
rect 3244 5958 3256 6010
rect 3308 5958 3320 6010
rect 3372 5958 3384 6010
rect 3436 5958 3448 6010
rect 3500 5958 4687 6010
rect 4739 5958 4751 6010
rect 4803 5958 4815 6010
rect 4867 5958 4879 6010
rect 4931 5958 4943 6010
rect 4995 5958 6182 6010
rect 6234 5958 6246 6010
rect 6298 5958 6310 6010
rect 6362 5958 6374 6010
rect 6426 5958 6438 6010
rect 6490 5958 7084 6010
rect 1104 5936 7084 5958
rect 5064 5899 5122 5905
rect 5064 5865 5076 5899
rect 5110 5896 5122 5899
rect 5534 5896 5540 5908
rect 5110 5868 5540 5896
rect 5110 5865 5122 5868
rect 5064 5859 5122 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 6546 5856 6552 5908
rect 6604 5856 6610 5908
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5729 2007 5763
rect 1949 5723 2007 5729
rect 1964 5692 1992 5723
rect 2038 5720 2044 5772
rect 2096 5720 2102 5772
rect 3050 5720 3056 5772
rect 3108 5720 3114 5772
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5760 4859 5763
rect 5166 5760 5172 5772
rect 4847 5732 5172 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 3068 5692 3096 5720
rect 1964 5664 3096 5692
rect 2133 5627 2191 5633
rect 2133 5593 2145 5627
rect 2179 5624 2191 5627
rect 2774 5624 2780 5636
rect 2179 5596 2780 5624
rect 2179 5593 2191 5596
rect 2133 5587 2191 5593
rect 2774 5584 2780 5596
rect 2832 5584 2838 5636
rect 6086 5584 6092 5636
rect 6144 5584 6150 5636
rect 2222 5516 2228 5568
rect 2280 5556 2286 5568
rect 2501 5559 2559 5565
rect 2501 5556 2513 5559
rect 2280 5528 2513 5556
rect 2280 5516 2286 5528
rect 2501 5525 2513 5528
rect 2547 5525 2559 5559
rect 2501 5519 2559 5525
rect 1104 5466 7156 5488
rect 1104 5414 2357 5466
rect 2409 5414 2421 5466
rect 2473 5414 2485 5466
rect 2537 5414 2549 5466
rect 2601 5414 2613 5466
rect 2665 5414 3852 5466
rect 3904 5414 3916 5466
rect 3968 5414 3980 5466
rect 4032 5414 4044 5466
rect 4096 5414 4108 5466
rect 4160 5414 5347 5466
rect 5399 5414 5411 5466
rect 5463 5414 5475 5466
rect 5527 5414 5539 5466
rect 5591 5414 5603 5466
rect 5655 5414 6842 5466
rect 6894 5414 6906 5466
rect 6958 5414 6970 5466
rect 7022 5414 7034 5466
rect 7086 5414 7098 5466
rect 7150 5414 7156 5466
rect 1104 5392 7156 5414
rect 2958 5352 2964 5364
rect 1780 5324 2964 5352
rect 1780 5293 1808 5324
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5258 5352 5264 5364
rect 5123 5324 5264 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6086 5352 6092 5364
rect 6043 5324 6092 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5253 1823 5287
rect 3694 5284 3700 5296
rect 3542 5256 3700 5284
rect 1765 5247 1823 5253
rect 3694 5244 3700 5256
rect 3752 5244 3758 5296
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5132 5188 5457 5216
rect 5132 5176 5138 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 5537 5219 5595 5225
rect 5537 5185 5549 5219
rect 5583 5216 5595 5219
rect 6089 5219 6147 5225
rect 5583 5188 6040 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 6012 5160 6040 5188
rect 6089 5185 6101 5219
rect 6135 5185 6147 5219
rect 6089 5179 6147 5185
rect 2038 5108 2044 5160
rect 2096 5108 2102 5160
rect 2314 5108 2320 5160
rect 2372 5108 2378 5160
rect 3789 5151 3847 5157
rect 3789 5117 3801 5151
rect 3835 5148 3847 5151
rect 4893 5151 4951 5157
rect 4893 5148 4905 5151
rect 3835 5120 4905 5148
rect 3835 5117 3847 5120
rect 3789 5111 3847 5117
rect 4893 5117 4905 5120
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5675 5120 5856 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 4908 5080 4936 5111
rect 5828 5092 5856 5120
rect 5994 5108 6000 5160
rect 6052 5108 6058 5160
rect 5718 5080 5724 5092
rect 4908 5052 5724 5080
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 5810 5040 5816 5092
rect 5868 5040 5874 5092
rect 5902 5040 5908 5092
rect 5960 5080 5966 5092
rect 6104 5080 6132 5179
rect 5960 5052 6132 5080
rect 5960 5040 5966 5052
rect 934 4972 940 5024
rect 992 5012 998 5024
rect 1489 5015 1547 5021
rect 1489 5012 1501 5015
rect 992 4984 1501 5012
rect 992 4972 998 4984
rect 1489 4981 1501 4984
rect 1535 4981 1547 5015
rect 1489 4975 1547 4981
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 6086 5012 6092 5024
rect 4387 4984 6092 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 1104 4922 7084 4944
rect 1104 4870 1697 4922
rect 1749 4870 1761 4922
rect 1813 4870 1825 4922
rect 1877 4870 1889 4922
rect 1941 4870 1953 4922
rect 2005 4870 3192 4922
rect 3244 4870 3256 4922
rect 3308 4870 3320 4922
rect 3372 4870 3384 4922
rect 3436 4870 3448 4922
rect 3500 4870 4687 4922
rect 4739 4870 4751 4922
rect 4803 4870 4815 4922
rect 4867 4870 4879 4922
rect 4931 4870 4943 4922
rect 4995 4870 6182 4922
rect 6234 4870 6246 4922
rect 6298 4870 6310 4922
rect 6362 4870 6374 4922
rect 6426 4870 6438 4922
rect 6490 4870 7084 4922
rect 1104 4848 7084 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2314 4808 2320 4820
rect 1995 4780 2320 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2777 4743 2835 4749
rect 2777 4709 2789 4743
rect 2823 4709 2835 4743
rect 2777 4703 2835 4709
rect 2792 4672 2820 4703
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 5810 4740 5816 4752
rect 3108 4712 5816 4740
rect 3108 4700 3114 4712
rect 3436 4681 3464 4712
rect 5810 4700 5816 4712
rect 5868 4740 5874 4752
rect 5868 4712 6224 4740
rect 5868 4700 5874 4712
rect 1780 4644 2820 4672
rect 3421 4675 3479 4681
rect 1780 4613 1808 4644
rect 3421 4641 3433 4675
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 6086 4632 6092 4684
rect 6144 4632 6150 4684
rect 6196 4681 6224 4712
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4573 1823 4607
rect 1765 4567 1823 4573
rect 2222 4564 2228 4616
rect 2280 4564 2286 4616
rect 2774 4564 2780 4616
rect 2832 4604 2838 4616
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 2832 4576 3249 4604
rect 2832 4564 2838 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 3789 4539 3847 4545
rect 3789 4536 3801 4539
rect 2924 4508 3801 4536
rect 2924 4496 2930 4508
rect 3789 4505 3801 4508
rect 3835 4505 3847 4539
rect 6104 4536 6132 4632
rect 3789 4499 3847 4505
rect 4540 4508 6132 4536
rect 2041 4471 2099 4477
rect 2041 4437 2053 4471
rect 2087 4468 2099 4471
rect 2130 4468 2136 4480
rect 2087 4440 2136 4468
rect 2087 4437 2099 4440
rect 2041 4431 2099 4437
rect 2130 4428 2136 4440
rect 2188 4428 2194 4480
rect 3145 4471 3203 4477
rect 3145 4437 3157 4471
rect 3191 4468 3203 4471
rect 4540 4468 4568 4508
rect 3191 4440 4568 4468
rect 3191 4437 3203 4440
rect 3145 4431 3203 4437
rect 5074 4428 5080 4480
rect 5132 4428 5138 4480
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5629 4471 5687 4477
rect 5629 4468 5641 4471
rect 5316 4440 5641 4468
rect 5316 4428 5322 4440
rect 5629 4437 5641 4440
rect 5675 4437 5687 4471
rect 5629 4431 5687 4437
rect 5994 4428 6000 4480
rect 6052 4428 6058 4480
rect 1104 4378 7156 4400
rect 1104 4326 2357 4378
rect 2409 4326 2421 4378
rect 2473 4326 2485 4378
rect 2537 4326 2549 4378
rect 2601 4326 2613 4378
rect 2665 4326 3852 4378
rect 3904 4326 3916 4378
rect 3968 4326 3980 4378
rect 4032 4326 4044 4378
rect 4096 4326 4108 4378
rect 4160 4326 5347 4378
rect 5399 4326 5411 4378
rect 5463 4326 5475 4378
rect 5527 4326 5539 4378
rect 5591 4326 5603 4378
rect 5655 4326 6842 4378
rect 6894 4326 6906 4378
rect 6958 4326 6970 4378
rect 7022 4326 7034 4378
rect 7086 4326 7098 4378
rect 7150 4326 7156 4378
rect 1104 4304 7156 4326
rect 2774 4224 2780 4276
rect 2832 4224 2838 4276
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 3881 4267 3939 4273
rect 3881 4264 3893 4267
rect 3752 4236 3893 4264
rect 3752 4224 3758 4236
rect 3881 4233 3893 4236
rect 3927 4233 3939 4267
rect 3881 4227 3939 4233
rect 5718 4224 5724 4276
rect 5776 4224 5782 4276
rect 5736 4196 5764 4224
rect 5813 4199 5871 4205
rect 5813 4196 5825 4199
rect 5736 4168 5825 4196
rect 5813 4165 5825 4168
rect 5859 4165 5871 4199
rect 5813 4159 5871 4165
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3016 4100 3341 4128
rect 3016 4088 3022 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 3988 4060 4016 4091
rect 5810 4060 5816 4072
rect 3988 4032 5816 4060
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6089 4063 6147 4069
rect 6089 4029 6101 4063
rect 6135 4060 6147 4063
rect 7282 4060 7288 4072
rect 6135 4032 7288 4060
rect 6135 4029 6147 4032
rect 6089 4023 6147 4029
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 1104 3834 7084 3856
rect 1104 3782 1697 3834
rect 1749 3782 1761 3834
rect 1813 3782 1825 3834
rect 1877 3782 1889 3834
rect 1941 3782 1953 3834
rect 2005 3782 3192 3834
rect 3244 3782 3256 3834
rect 3308 3782 3320 3834
rect 3372 3782 3384 3834
rect 3436 3782 3448 3834
rect 3500 3782 4687 3834
rect 4739 3782 4751 3834
rect 4803 3782 4815 3834
rect 4867 3782 4879 3834
rect 4931 3782 4943 3834
rect 4995 3782 6182 3834
rect 6234 3782 6246 3834
rect 6298 3782 6310 3834
rect 6362 3782 6374 3834
rect 6426 3782 6438 3834
rect 6490 3782 7084 3834
rect 1104 3760 7084 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3016 3692 3433 3720
rect 3016 3680 3022 3692
rect 3421 3689 3433 3692
rect 3467 3689 3479 3723
rect 3421 3683 3479 3689
rect 5258 3680 5264 3732
rect 5316 3680 5322 3732
rect 1673 3587 1731 3593
rect 1673 3553 1685 3587
rect 1719 3584 1731 3587
rect 2038 3584 2044 3596
rect 1719 3556 2044 3584
rect 1719 3553 1731 3556
rect 1673 3547 1731 3553
rect 2038 3544 2044 3556
rect 2096 3544 2102 3596
rect 5276 3584 5304 3680
rect 4816 3556 5304 3584
rect 4816 3525 4844 3556
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3417 2007 3451
rect 3326 3448 3332 3460
rect 3174 3420 3332 3448
rect 1949 3411 2007 3417
rect 1964 3380 1992 3411
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 5276 3448 5304 3479
rect 5810 3448 5816 3460
rect 5276 3420 5816 3448
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 2130 3380 2136 3392
rect 1964 3352 2136 3380
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 4522 3340 4528 3392
rect 4580 3380 4586 3392
rect 4617 3383 4675 3389
rect 4617 3380 4629 3383
rect 4580 3352 4629 3380
rect 4580 3340 4586 3352
rect 4617 3349 4629 3352
rect 4663 3349 4675 3383
rect 4617 3343 4675 3349
rect 5353 3383 5411 3389
rect 5353 3349 5365 3383
rect 5399 3380 5411 3383
rect 5718 3380 5724 3392
rect 5399 3352 5724 3380
rect 5399 3349 5411 3352
rect 5353 3343 5411 3349
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 1104 3290 7156 3312
rect 1104 3238 2357 3290
rect 2409 3238 2421 3290
rect 2473 3238 2485 3290
rect 2537 3238 2549 3290
rect 2601 3238 2613 3290
rect 2665 3238 3852 3290
rect 3904 3238 3916 3290
rect 3968 3238 3980 3290
rect 4032 3238 4044 3290
rect 4096 3238 4108 3290
rect 4160 3238 5347 3290
rect 5399 3238 5411 3290
rect 5463 3238 5475 3290
rect 5527 3238 5539 3290
rect 5591 3238 5603 3290
rect 5655 3238 6842 3290
rect 6894 3238 6906 3290
rect 6958 3238 6970 3290
rect 7022 3238 7034 3290
rect 7086 3238 7098 3290
rect 7150 3238 7156 3290
rect 1104 3216 7156 3238
rect 1857 3179 1915 3185
rect 1857 3145 1869 3179
rect 1903 3176 1915 3179
rect 2038 3176 2044 3188
rect 1903 3148 2044 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 3326 3136 3332 3188
rect 3384 3136 3390 3188
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 5224 3148 5733 3176
rect 5224 3136 5230 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 3145 3111 3203 3117
rect 3145 3077 3157 3111
rect 3191 3108 3203 3111
rect 4433 3111 4491 3117
rect 4433 3108 4445 3111
rect 3191 3080 4445 3108
rect 3191 3077 3203 3080
rect 3145 3071 3203 3077
rect 4433 3077 4445 3080
rect 4479 3108 4491 3111
rect 5074 3108 5080 3120
rect 4479 3080 5080 3108
rect 4479 3077 4491 3080
rect 4433 3071 4491 3077
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3421 3003 3479 3009
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 3436 2904 3464 3003
rect 4080 2972 4108 3003
rect 5994 2972 6000 2984
rect 4080 2944 6000 2972
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 5810 2904 5816 2916
rect 3436 2876 5816 2904
rect 5810 2864 5816 2876
rect 5868 2864 5874 2916
rect 3973 2839 4031 2845
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 4338 2836 4344 2848
rect 4019 2808 4344 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 1104 2746 7084 2768
rect 1104 2694 1697 2746
rect 1749 2694 1761 2746
rect 1813 2694 1825 2746
rect 1877 2694 1889 2746
rect 1941 2694 1953 2746
rect 2005 2694 3192 2746
rect 3244 2694 3256 2746
rect 3308 2694 3320 2746
rect 3372 2694 3384 2746
rect 3436 2694 3448 2746
rect 3500 2694 4687 2746
rect 4739 2694 4751 2746
rect 4803 2694 4815 2746
rect 4867 2694 4879 2746
rect 4931 2694 4943 2746
rect 4995 2694 6182 2746
rect 6234 2694 6246 2746
rect 6298 2694 6310 2746
rect 6362 2694 6374 2746
rect 6426 2694 6438 2746
rect 6490 2694 7084 2746
rect 1104 2672 7084 2694
rect 5994 2592 6000 2644
rect 6052 2592 6058 2644
rect 5810 2524 5816 2576
rect 5868 2564 5874 2576
rect 6457 2567 6515 2573
rect 6457 2564 6469 2567
rect 5868 2536 6469 2564
rect 5868 2524 5874 2536
rect 6457 2533 6469 2536
rect 6503 2533 6515 2567
rect 6457 2527 6515 2533
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 5166 2496 5172 2508
rect 4295 2468 5172 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5718 2456 5724 2508
rect 5776 2456 5782 2508
rect 5736 2428 5764 2456
rect 5658 2400 5764 2428
rect 4522 2320 4528 2372
rect 4580 2320 4586 2372
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 7190 2360 7196 2372
rect 6687 2332 7196 2360
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 1104 2202 7156 2224
rect 1104 2150 2357 2202
rect 2409 2150 2421 2202
rect 2473 2150 2485 2202
rect 2537 2150 2549 2202
rect 2601 2150 2613 2202
rect 2665 2150 3852 2202
rect 3904 2150 3916 2202
rect 3968 2150 3980 2202
rect 4032 2150 4044 2202
rect 4096 2150 4108 2202
rect 4160 2150 5347 2202
rect 5399 2150 5411 2202
rect 5463 2150 5475 2202
rect 5527 2150 5539 2202
rect 5591 2150 5603 2202
rect 5655 2150 6842 2202
rect 6894 2150 6906 2202
rect 6958 2150 6970 2202
rect 7022 2150 7034 2202
rect 7086 2150 7098 2202
rect 7150 2150 7156 2202
rect 1104 2128 7156 2150
<< via1 >>
rect 1697 8134 1749 8186
rect 1761 8134 1813 8186
rect 1825 8134 1877 8186
rect 1889 8134 1941 8186
rect 1953 8134 2005 8186
rect 3192 8134 3244 8186
rect 3256 8134 3308 8186
rect 3320 8134 3372 8186
rect 3384 8134 3436 8186
rect 3448 8134 3500 8186
rect 4687 8134 4739 8186
rect 4751 8134 4803 8186
rect 4815 8134 4867 8186
rect 4879 8134 4931 8186
rect 4943 8134 4995 8186
rect 6182 8134 6234 8186
rect 6246 8134 6298 8186
rect 6310 8134 6362 8186
rect 6374 8134 6426 8186
rect 6438 8134 6490 8186
rect 7748 8032 7800 8084
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 3608 7828 3660 7880
rect 6092 7803 6144 7812
rect 6092 7769 6101 7803
rect 6101 7769 6135 7803
rect 6135 7769 6144 7803
rect 6092 7760 6144 7769
rect 2044 7692 2096 7744
rect 3056 7692 3108 7744
rect 2357 7590 2409 7642
rect 2421 7590 2473 7642
rect 2485 7590 2537 7642
rect 2549 7590 2601 7642
rect 2613 7590 2665 7642
rect 3852 7590 3904 7642
rect 3916 7590 3968 7642
rect 3980 7590 4032 7642
rect 4044 7590 4096 7642
rect 4108 7590 4160 7642
rect 5347 7590 5399 7642
rect 5411 7590 5463 7642
rect 5475 7590 5527 7642
rect 5539 7590 5591 7642
rect 5603 7590 5655 7642
rect 6842 7590 6894 7642
rect 6906 7590 6958 7642
rect 6970 7590 7022 7642
rect 7034 7590 7086 7642
rect 7098 7590 7150 7642
rect 1697 7046 1749 7098
rect 1761 7046 1813 7098
rect 1825 7046 1877 7098
rect 1889 7046 1941 7098
rect 1953 7046 2005 7098
rect 3192 7046 3244 7098
rect 3256 7046 3308 7098
rect 3320 7046 3372 7098
rect 3384 7046 3436 7098
rect 3448 7046 3500 7098
rect 4687 7046 4739 7098
rect 4751 7046 4803 7098
rect 4815 7046 4867 7098
rect 4879 7046 4931 7098
rect 4943 7046 4995 7098
rect 6182 7046 6234 7098
rect 6246 7046 6298 7098
rect 6310 7046 6362 7098
rect 6374 7046 6426 7098
rect 6438 7046 6490 7098
rect 6092 6808 6144 6860
rect 6552 6808 6604 6860
rect 5080 6604 5132 6656
rect 2357 6502 2409 6554
rect 2421 6502 2473 6554
rect 2485 6502 2537 6554
rect 2549 6502 2601 6554
rect 2613 6502 2665 6554
rect 3852 6502 3904 6554
rect 3916 6502 3968 6554
rect 3980 6502 4032 6554
rect 4044 6502 4096 6554
rect 4108 6502 4160 6554
rect 5347 6502 5399 6554
rect 5411 6502 5463 6554
rect 5475 6502 5527 6554
rect 5539 6502 5591 6554
rect 5603 6502 5655 6554
rect 6842 6502 6894 6554
rect 6906 6502 6958 6554
rect 6970 6502 7022 6554
rect 7034 6502 7086 6554
rect 7098 6502 7150 6554
rect 5264 6239 5316 6248
rect 5264 6205 5273 6239
rect 5273 6205 5307 6239
rect 5307 6205 5316 6239
rect 5264 6196 5316 6205
rect 5540 6060 5592 6112
rect 1697 5958 1749 6010
rect 1761 5958 1813 6010
rect 1825 5958 1877 6010
rect 1889 5958 1941 6010
rect 1953 5958 2005 6010
rect 3192 5958 3244 6010
rect 3256 5958 3308 6010
rect 3320 5958 3372 6010
rect 3384 5958 3436 6010
rect 3448 5958 3500 6010
rect 4687 5958 4739 6010
rect 4751 5958 4803 6010
rect 4815 5958 4867 6010
rect 4879 5958 4931 6010
rect 4943 5958 4995 6010
rect 6182 5958 6234 6010
rect 6246 5958 6298 6010
rect 6310 5958 6362 6010
rect 6374 5958 6426 6010
rect 6438 5958 6490 6010
rect 5540 5856 5592 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 2044 5763 2096 5772
rect 2044 5729 2053 5763
rect 2053 5729 2087 5763
rect 2087 5729 2096 5763
rect 2044 5720 2096 5729
rect 3056 5720 3108 5772
rect 5172 5720 5224 5772
rect 2780 5584 2832 5636
rect 6092 5584 6144 5636
rect 2228 5516 2280 5568
rect 2357 5414 2409 5466
rect 2421 5414 2473 5466
rect 2485 5414 2537 5466
rect 2549 5414 2601 5466
rect 2613 5414 2665 5466
rect 3852 5414 3904 5466
rect 3916 5414 3968 5466
rect 3980 5414 4032 5466
rect 4044 5414 4096 5466
rect 4108 5414 4160 5466
rect 5347 5414 5399 5466
rect 5411 5414 5463 5466
rect 5475 5414 5527 5466
rect 5539 5414 5591 5466
rect 5603 5414 5655 5466
rect 6842 5414 6894 5466
rect 6906 5414 6958 5466
rect 6970 5414 7022 5466
rect 7034 5414 7086 5466
rect 7098 5414 7150 5466
rect 2964 5312 3016 5364
rect 5264 5312 5316 5364
rect 6092 5312 6144 5364
rect 3700 5244 3752 5296
rect 5080 5176 5132 5228
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 2320 5151 2372 5160
rect 2320 5117 2329 5151
rect 2329 5117 2363 5151
rect 2363 5117 2372 5151
rect 2320 5108 2372 5117
rect 6000 5108 6052 5160
rect 5724 5040 5776 5092
rect 5816 5040 5868 5092
rect 5908 5040 5960 5092
rect 940 4972 992 5024
rect 6092 4972 6144 5024
rect 1697 4870 1749 4922
rect 1761 4870 1813 4922
rect 1825 4870 1877 4922
rect 1889 4870 1941 4922
rect 1953 4870 2005 4922
rect 3192 4870 3244 4922
rect 3256 4870 3308 4922
rect 3320 4870 3372 4922
rect 3384 4870 3436 4922
rect 3448 4870 3500 4922
rect 4687 4870 4739 4922
rect 4751 4870 4803 4922
rect 4815 4870 4867 4922
rect 4879 4870 4931 4922
rect 4943 4870 4995 4922
rect 6182 4870 6234 4922
rect 6246 4870 6298 4922
rect 6310 4870 6362 4922
rect 6374 4870 6426 4922
rect 6438 4870 6490 4922
rect 2320 4768 2372 4820
rect 3056 4700 3108 4752
rect 5816 4700 5868 4752
rect 6092 4675 6144 4684
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 2780 4564 2832 4616
rect 2872 4496 2924 4548
rect 2136 4428 2188 4480
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 5264 4428 5316 4480
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 2357 4326 2409 4378
rect 2421 4326 2473 4378
rect 2485 4326 2537 4378
rect 2549 4326 2601 4378
rect 2613 4326 2665 4378
rect 3852 4326 3904 4378
rect 3916 4326 3968 4378
rect 3980 4326 4032 4378
rect 4044 4326 4096 4378
rect 4108 4326 4160 4378
rect 5347 4326 5399 4378
rect 5411 4326 5463 4378
rect 5475 4326 5527 4378
rect 5539 4326 5591 4378
rect 5603 4326 5655 4378
rect 6842 4326 6894 4378
rect 6906 4326 6958 4378
rect 6970 4326 7022 4378
rect 7034 4326 7086 4378
rect 7098 4326 7150 4378
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 3700 4224 3752 4276
rect 5724 4224 5776 4276
rect 2964 4088 3016 4140
rect 5816 4020 5868 4072
rect 7288 4020 7340 4072
rect 1697 3782 1749 3834
rect 1761 3782 1813 3834
rect 1825 3782 1877 3834
rect 1889 3782 1941 3834
rect 1953 3782 2005 3834
rect 3192 3782 3244 3834
rect 3256 3782 3308 3834
rect 3320 3782 3372 3834
rect 3384 3782 3436 3834
rect 3448 3782 3500 3834
rect 4687 3782 4739 3834
rect 4751 3782 4803 3834
rect 4815 3782 4867 3834
rect 4879 3782 4931 3834
rect 4943 3782 4995 3834
rect 6182 3782 6234 3834
rect 6246 3782 6298 3834
rect 6310 3782 6362 3834
rect 6374 3782 6426 3834
rect 6438 3782 6490 3834
rect 2964 3680 3016 3732
rect 5264 3680 5316 3732
rect 2044 3544 2096 3596
rect 3332 3408 3384 3460
rect 5816 3408 5868 3460
rect 2136 3340 2188 3392
rect 4528 3340 4580 3392
rect 5724 3340 5776 3392
rect 2357 3238 2409 3290
rect 2421 3238 2473 3290
rect 2485 3238 2537 3290
rect 2549 3238 2601 3290
rect 2613 3238 2665 3290
rect 3852 3238 3904 3290
rect 3916 3238 3968 3290
rect 3980 3238 4032 3290
rect 4044 3238 4096 3290
rect 4108 3238 4160 3290
rect 5347 3238 5399 3290
rect 5411 3238 5463 3290
rect 5475 3238 5527 3290
rect 5539 3238 5591 3290
rect 5603 3238 5655 3290
rect 6842 3238 6894 3290
rect 6906 3238 6958 3290
rect 6970 3238 7022 3290
rect 7034 3238 7086 3290
rect 7098 3238 7150 3290
rect 2044 3136 2096 3188
rect 3332 3179 3384 3188
rect 3332 3145 3341 3179
rect 3341 3145 3375 3179
rect 3375 3145 3384 3179
rect 3332 3136 3384 3145
rect 5172 3136 5224 3188
rect 5080 3068 5132 3120
rect 6000 2932 6052 2984
rect 5816 2864 5868 2916
rect 4344 2796 4396 2848
rect 1697 2694 1749 2746
rect 1761 2694 1813 2746
rect 1825 2694 1877 2746
rect 1889 2694 1941 2746
rect 1953 2694 2005 2746
rect 3192 2694 3244 2746
rect 3256 2694 3308 2746
rect 3320 2694 3372 2746
rect 3384 2694 3436 2746
rect 3448 2694 3500 2746
rect 4687 2694 4739 2746
rect 4751 2694 4803 2746
rect 4815 2694 4867 2746
rect 4879 2694 4931 2746
rect 4943 2694 4995 2746
rect 6182 2694 6234 2746
rect 6246 2694 6298 2746
rect 6310 2694 6362 2746
rect 6374 2694 6426 2746
rect 6438 2694 6490 2746
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 5816 2524 5868 2576
rect 5172 2456 5224 2508
rect 5724 2456 5776 2508
rect 4528 2363 4580 2372
rect 4528 2329 4537 2363
rect 4537 2329 4571 2363
rect 4571 2329 4580 2363
rect 4528 2320 4580 2329
rect 7196 2320 7248 2372
rect 2357 2150 2409 2202
rect 2421 2150 2473 2202
rect 2485 2150 2537 2202
rect 2549 2150 2601 2202
rect 2613 2150 2665 2202
rect 3852 2150 3904 2202
rect 3916 2150 3968 2202
rect 3980 2150 4032 2202
rect 4044 2150 4096 2202
rect 4108 2150 4160 2202
rect 5347 2150 5399 2202
rect 5411 2150 5463 2202
rect 5475 2150 5527 2202
rect 5539 2150 5591 2202
rect 5603 2150 5655 2202
rect 6842 2150 6894 2202
rect 6906 2150 6958 2202
rect 6970 2150 7022 2202
rect 7034 2150 7086 2202
rect 7098 2150 7150 2202
<< metal2 >>
rect 3238 9555 3294 10355
rect 3344 9574 3648 9602
rect 1398 9480 1454 9489
rect 3252 9466 3280 9555
rect 3344 9466 3372 9574
rect 3252 9438 3372 9466
rect 1398 9415 1454 9424
rect 1412 7886 1440 9415
rect 1697 8188 2005 8197
rect 1697 8186 1703 8188
rect 1759 8186 1783 8188
rect 1839 8186 1863 8188
rect 1919 8186 1943 8188
rect 1999 8186 2005 8188
rect 1759 8134 1761 8186
rect 1941 8134 1943 8186
rect 1697 8132 1703 8134
rect 1759 8132 1783 8134
rect 1839 8132 1863 8134
rect 1919 8132 1943 8134
rect 1999 8132 2005 8134
rect 1697 8123 2005 8132
rect 3192 8188 3500 8197
rect 3192 8186 3198 8188
rect 3254 8186 3278 8188
rect 3334 8186 3358 8188
rect 3414 8186 3438 8188
rect 3494 8186 3500 8188
rect 3254 8134 3256 8186
rect 3436 8134 3438 8186
rect 3192 8132 3198 8134
rect 3254 8132 3278 8134
rect 3334 8132 3358 8134
rect 3414 8132 3438 8134
rect 3494 8132 3500 8134
rect 3192 8123 3500 8132
rect 3620 7886 3648 9574
rect 7746 9555 7802 10355
rect 4687 8188 4995 8197
rect 4687 8186 4693 8188
rect 4749 8186 4773 8188
rect 4829 8186 4853 8188
rect 4909 8186 4933 8188
rect 4989 8186 4995 8188
rect 4749 8134 4751 8186
rect 4931 8134 4933 8186
rect 4687 8132 4693 8134
rect 4749 8132 4773 8134
rect 4829 8132 4853 8134
rect 4909 8132 4933 8134
rect 4989 8132 4995 8134
rect 4687 8123 4995 8132
rect 6182 8188 6490 8197
rect 6182 8186 6188 8188
rect 6244 8186 6268 8188
rect 6324 8186 6348 8188
rect 6404 8186 6428 8188
rect 6484 8186 6490 8188
rect 6244 8134 6246 8186
rect 6426 8134 6428 8186
rect 6182 8132 6188 8134
rect 6244 8132 6268 8134
rect 6324 8132 6348 8134
rect 6404 8132 6428 8134
rect 6484 8132 6490 8134
rect 6182 8123 6490 8132
rect 7760 8090 7788 9555
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 3056 7744 3108 7750
rect 3056 7686 3108 7692
rect 1697 7100 2005 7109
rect 1697 7098 1703 7100
rect 1759 7098 1783 7100
rect 1839 7098 1863 7100
rect 1919 7098 1943 7100
rect 1999 7098 2005 7100
rect 1759 7046 1761 7098
rect 1941 7046 1943 7098
rect 1697 7044 1703 7046
rect 1759 7044 1783 7046
rect 1839 7044 1863 7046
rect 1919 7044 1943 7046
rect 1999 7044 2005 7046
rect 1697 7035 2005 7044
rect 1697 6012 2005 6021
rect 1697 6010 1703 6012
rect 1759 6010 1783 6012
rect 1839 6010 1863 6012
rect 1919 6010 1943 6012
rect 1999 6010 2005 6012
rect 1759 5958 1761 6010
rect 1941 5958 1943 6010
rect 1697 5956 1703 5958
rect 1759 5956 1783 5958
rect 1839 5956 1863 5958
rect 1919 5956 1943 5958
rect 1999 5956 2005 5958
rect 1697 5947 2005 5956
rect 2056 5778 2084 7686
rect 2357 7644 2665 7653
rect 2357 7642 2363 7644
rect 2419 7642 2443 7644
rect 2499 7642 2523 7644
rect 2579 7642 2603 7644
rect 2659 7642 2665 7644
rect 2419 7590 2421 7642
rect 2601 7590 2603 7642
rect 2357 7588 2363 7590
rect 2419 7588 2443 7590
rect 2499 7588 2523 7590
rect 2579 7588 2603 7590
rect 2659 7588 2665 7590
rect 2357 7579 2665 7588
rect 2357 6556 2665 6565
rect 2357 6554 2363 6556
rect 2419 6554 2443 6556
rect 2499 6554 2523 6556
rect 2579 6554 2603 6556
rect 2659 6554 2665 6556
rect 2419 6502 2421 6554
rect 2601 6502 2603 6554
rect 2357 6500 2363 6502
rect 2419 6500 2443 6502
rect 2499 6500 2523 6502
rect 2579 6500 2603 6502
rect 2659 6500 2665 6502
rect 2357 6491 2665 6500
rect 3068 5778 3096 7686
rect 3852 7644 4160 7653
rect 3852 7642 3858 7644
rect 3914 7642 3938 7644
rect 3994 7642 4018 7644
rect 4074 7642 4098 7644
rect 4154 7642 4160 7644
rect 3914 7590 3916 7642
rect 4096 7590 4098 7642
rect 3852 7588 3858 7590
rect 3914 7588 3938 7590
rect 3994 7588 4018 7590
rect 4074 7588 4098 7590
rect 4154 7588 4160 7590
rect 3852 7579 4160 7588
rect 5347 7644 5655 7653
rect 5347 7642 5353 7644
rect 5409 7642 5433 7644
rect 5489 7642 5513 7644
rect 5569 7642 5593 7644
rect 5649 7642 5655 7644
rect 5409 7590 5411 7642
rect 5591 7590 5593 7642
rect 5347 7588 5353 7590
rect 5409 7588 5433 7590
rect 5489 7588 5513 7590
rect 5569 7588 5593 7590
rect 5649 7588 5655 7590
rect 5347 7579 5655 7588
rect 3192 7100 3500 7109
rect 3192 7098 3198 7100
rect 3254 7098 3278 7100
rect 3334 7098 3358 7100
rect 3414 7098 3438 7100
rect 3494 7098 3500 7100
rect 3254 7046 3256 7098
rect 3436 7046 3438 7098
rect 3192 7044 3198 7046
rect 3254 7044 3278 7046
rect 3334 7044 3358 7046
rect 3414 7044 3438 7046
rect 3494 7044 3500 7046
rect 3192 7035 3500 7044
rect 4687 7100 4995 7109
rect 4687 7098 4693 7100
rect 4749 7098 4773 7100
rect 4829 7098 4853 7100
rect 4909 7098 4933 7100
rect 4989 7098 4995 7100
rect 4749 7046 4751 7098
rect 4931 7046 4933 7098
rect 4687 7044 4693 7046
rect 4749 7044 4773 7046
rect 4829 7044 4853 7046
rect 4909 7044 4933 7046
rect 4989 7044 4995 7046
rect 4687 7035 4995 7044
rect 6104 6866 6132 7754
rect 6842 7644 7150 7653
rect 6842 7642 6848 7644
rect 6904 7642 6928 7644
rect 6984 7642 7008 7644
rect 7064 7642 7088 7644
rect 7144 7642 7150 7644
rect 6904 7590 6906 7642
rect 7086 7590 7088 7642
rect 6842 7588 6848 7590
rect 6904 7588 6928 7590
rect 6984 7588 7008 7590
rect 7064 7588 7088 7590
rect 7144 7588 7150 7590
rect 6842 7579 7150 7588
rect 6182 7100 6490 7109
rect 6182 7098 6188 7100
rect 6244 7098 6268 7100
rect 6324 7098 6348 7100
rect 6404 7098 6428 7100
rect 6484 7098 6490 7100
rect 6244 7046 6246 7098
rect 6426 7046 6428 7098
rect 6182 7044 6188 7046
rect 6244 7044 6268 7046
rect 6324 7044 6348 7046
rect 6404 7044 6428 7046
rect 6484 7044 6490 7046
rect 6182 7035 6490 7044
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 3852 6556 4160 6565
rect 3852 6554 3858 6556
rect 3914 6554 3938 6556
rect 3994 6554 4018 6556
rect 4074 6554 4098 6556
rect 4154 6554 4160 6556
rect 3914 6502 3916 6554
rect 4096 6502 4098 6554
rect 3852 6500 3858 6502
rect 3914 6500 3938 6502
rect 3994 6500 4018 6502
rect 4074 6500 4098 6502
rect 4154 6500 4160 6502
rect 3852 6491 4160 6500
rect 3192 6012 3500 6021
rect 3192 6010 3198 6012
rect 3254 6010 3278 6012
rect 3334 6010 3358 6012
rect 3414 6010 3438 6012
rect 3494 6010 3500 6012
rect 3254 5958 3256 6010
rect 3436 5958 3438 6010
rect 3192 5956 3198 5958
rect 3254 5956 3278 5958
rect 3334 5956 3358 5958
rect 3414 5956 3438 5958
rect 3494 5956 3500 5958
rect 3192 5947 3500 5956
rect 4687 6012 4995 6021
rect 4687 6010 4693 6012
rect 4749 6010 4773 6012
rect 4829 6010 4853 6012
rect 4909 6010 4933 6012
rect 4989 6010 4995 6012
rect 4749 5958 4751 6010
rect 4931 5958 4933 6010
rect 4687 5956 4693 5958
rect 4749 5956 4773 5958
rect 4829 5956 4853 5958
rect 4909 5956 4933 5958
rect 4989 5956 4995 5958
rect 4687 5947 4995 5956
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 940 5024 992 5030
rect 940 4966 992 4972
rect 952 4865 980 4966
rect 1697 4924 2005 4933
rect 1697 4922 1703 4924
rect 1759 4922 1783 4924
rect 1839 4922 1863 4924
rect 1919 4922 1943 4924
rect 1999 4922 2005 4924
rect 1759 4870 1761 4922
rect 1941 4870 1943 4922
rect 1697 4868 1703 4870
rect 1759 4868 1783 4870
rect 1839 4868 1863 4870
rect 1919 4868 1943 4870
rect 1999 4868 2005 4870
rect 938 4856 994 4865
rect 1697 4859 2005 4868
rect 938 4791 994 4800
rect 1697 3836 2005 3845
rect 1697 3834 1703 3836
rect 1759 3834 1783 3836
rect 1839 3834 1863 3836
rect 1919 3834 1943 3836
rect 1999 3834 2005 3836
rect 1759 3782 1761 3834
rect 1941 3782 1943 3834
rect 1697 3780 1703 3782
rect 1759 3780 1783 3782
rect 1839 3780 1863 3782
rect 1919 3780 1943 3782
rect 1999 3780 2005 3782
rect 1697 3771 2005 3780
rect 2056 3602 2084 5102
rect 2240 4622 2268 5510
rect 2357 5468 2665 5477
rect 2357 5466 2363 5468
rect 2419 5466 2443 5468
rect 2499 5466 2523 5468
rect 2579 5466 2603 5468
rect 2659 5466 2665 5468
rect 2419 5414 2421 5466
rect 2601 5414 2603 5466
rect 2357 5412 2363 5414
rect 2419 5412 2443 5414
rect 2499 5412 2523 5414
rect 2579 5412 2603 5414
rect 2659 5412 2665 5414
rect 2357 5403 2665 5412
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2332 4826 2360 5102
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2792 4622 2820 5578
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 2056 3194 2084 3538
rect 2148 3398 2176 4422
rect 2357 4380 2665 4389
rect 2357 4378 2363 4380
rect 2419 4378 2443 4380
rect 2499 4378 2523 4380
rect 2579 4378 2603 4380
rect 2659 4378 2665 4380
rect 2419 4326 2421 4378
rect 2601 4326 2603 4378
rect 2357 4324 2363 4326
rect 2419 4324 2443 4326
rect 2499 4324 2523 4326
rect 2579 4324 2603 4326
rect 2659 4324 2665 4326
rect 2357 4315 2665 4324
rect 2792 4282 2820 4558
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2357 3292 2665 3301
rect 2357 3290 2363 3292
rect 2419 3290 2443 3292
rect 2499 3290 2523 3292
rect 2579 3290 2603 3292
rect 2659 3290 2665 3292
rect 2419 3238 2421 3290
rect 2601 3238 2603 3290
rect 2357 3236 2363 3238
rect 2419 3236 2443 3238
rect 2499 3236 2523 3238
rect 2579 3236 2603 3238
rect 2659 3236 2665 3238
rect 2357 3227 2665 3236
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2884 2961 2912 4490
rect 2976 4146 3004 5306
rect 3068 4758 3096 5714
rect 3852 5468 4160 5477
rect 3852 5466 3858 5468
rect 3914 5466 3938 5468
rect 3994 5466 4018 5468
rect 4074 5466 4098 5468
rect 4154 5466 4160 5468
rect 3914 5414 3916 5466
rect 4096 5414 4098 5466
rect 3852 5412 3858 5414
rect 3914 5412 3938 5414
rect 3994 5412 4018 5414
rect 4074 5412 4098 5414
rect 4154 5412 4160 5414
rect 3852 5403 4160 5412
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3192 4924 3500 4933
rect 3192 4922 3198 4924
rect 3254 4922 3278 4924
rect 3334 4922 3358 4924
rect 3414 4922 3438 4924
rect 3494 4922 3500 4924
rect 3254 4870 3256 4922
rect 3436 4870 3438 4922
rect 3192 4868 3198 4870
rect 3254 4868 3278 4870
rect 3334 4868 3358 4870
rect 3414 4868 3438 4870
rect 3494 4868 3500 4870
rect 3192 4859 3500 4868
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3712 4282 3740 5238
rect 5092 5234 5120 6598
rect 5347 6556 5655 6565
rect 5347 6554 5353 6556
rect 5409 6554 5433 6556
rect 5489 6554 5513 6556
rect 5569 6554 5593 6556
rect 5649 6554 5655 6556
rect 5409 6502 5411 6554
rect 5591 6502 5593 6554
rect 5347 6500 5353 6502
rect 5409 6500 5433 6502
rect 5489 6500 5513 6502
rect 5569 6500 5593 6502
rect 5649 6500 5655 6502
rect 5347 6491 5655 6500
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4687 4924 4995 4933
rect 4687 4922 4693 4924
rect 4749 4922 4773 4924
rect 4829 4922 4853 4924
rect 4909 4922 4933 4924
rect 4989 4922 4995 4924
rect 4749 4870 4751 4922
rect 4931 4870 4933 4922
rect 4687 4868 4693 4870
rect 4749 4868 4773 4870
rect 4829 4868 4853 4870
rect 4909 4868 4933 4870
rect 4989 4868 4995 4870
rect 4687 4859 4995 4868
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 3852 4380 4160 4389
rect 3852 4378 3858 4380
rect 3914 4378 3938 4380
rect 3994 4378 4018 4380
rect 4074 4378 4098 4380
rect 4154 4378 4160 4380
rect 3914 4326 3916 4378
rect 4096 4326 4098 4378
rect 3852 4324 3858 4326
rect 3914 4324 3938 4326
rect 3994 4324 4018 4326
rect 4074 4324 4098 4326
rect 4154 4324 4160 4326
rect 3852 4315 4160 4324
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2976 3738 3004 4082
rect 3192 3836 3500 3845
rect 3192 3834 3198 3836
rect 3254 3834 3278 3836
rect 3334 3834 3358 3836
rect 3414 3834 3438 3836
rect 3494 3834 3500 3836
rect 3254 3782 3256 3834
rect 3436 3782 3438 3834
rect 3192 3780 3198 3782
rect 3254 3780 3278 3782
rect 3334 3780 3358 3782
rect 3414 3780 3438 3782
rect 3494 3780 3500 3782
rect 3192 3771 3500 3780
rect 4687 3836 4995 3845
rect 4687 3834 4693 3836
rect 4749 3834 4773 3836
rect 4829 3834 4853 3836
rect 4909 3834 4933 3836
rect 4989 3834 4995 3836
rect 4749 3782 4751 3834
rect 4931 3782 4933 3834
rect 4687 3780 4693 3782
rect 4749 3780 4773 3782
rect 4829 3780 4853 3782
rect 4909 3780 4933 3782
rect 4989 3780 4995 3782
rect 4687 3771 4995 3780
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3344 3194 3372 3402
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 3852 3292 4160 3301
rect 3852 3290 3858 3292
rect 3914 3290 3938 3292
rect 3994 3290 4018 3292
rect 4074 3290 4098 3292
rect 4154 3290 4160 3292
rect 3914 3238 3916 3290
rect 4096 3238 4098 3290
rect 3852 3236 3858 3238
rect 3914 3236 3938 3238
rect 3994 3236 4018 3238
rect 4074 3236 4098 3238
rect 4154 3236 4160 3238
rect 3852 3227 4160 3236
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 18 2952 74 2961
rect 18 2887 74 2896
rect 2870 2952 2926 2961
rect 2870 2887 2926 2896
rect 32 800 60 2887
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 1697 2748 2005 2757
rect 1697 2746 1703 2748
rect 1759 2746 1783 2748
rect 1839 2746 1863 2748
rect 1919 2746 1943 2748
rect 1999 2746 2005 2748
rect 1759 2694 1761 2746
rect 1941 2694 1943 2746
rect 1697 2692 1703 2694
rect 1759 2692 1783 2694
rect 1839 2692 1863 2694
rect 1919 2692 1943 2694
rect 1999 2692 2005 2694
rect 1697 2683 2005 2692
rect 3192 2748 3500 2757
rect 3192 2746 3198 2748
rect 3254 2746 3278 2748
rect 3334 2746 3358 2748
rect 3414 2746 3438 2748
rect 3494 2746 3500 2748
rect 3254 2694 3256 2746
rect 3436 2694 3438 2746
rect 3192 2692 3198 2694
rect 3254 2692 3278 2694
rect 3334 2692 3358 2694
rect 3414 2692 3438 2694
rect 3494 2692 3500 2694
rect 3192 2683 3500 2692
rect 2357 2204 2665 2213
rect 2357 2202 2363 2204
rect 2419 2202 2443 2204
rect 2499 2202 2523 2204
rect 2579 2202 2603 2204
rect 2659 2202 2665 2204
rect 2419 2150 2421 2202
rect 2601 2150 2603 2202
rect 2357 2148 2363 2150
rect 2419 2148 2443 2150
rect 2499 2148 2523 2150
rect 2579 2148 2603 2150
rect 2659 2148 2665 2150
rect 2357 2139 2665 2148
rect 3852 2204 4160 2213
rect 3852 2202 3858 2204
rect 3914 2202 3938 2204
rect 3994 2202 4018 2204
rect 4074 2202 4098 2204
rect 4154 2202 4160 2204
rect 3914 2150 3916 2202
rect 4096 2150 4098 2202
rect 3852 2148 3858 2150
rect 3914 2148 3938 2150
rect 3994 2148 4018 2150
rect 4074 2148 4098 2150
rect 4154 2148 4160 2150
rect 3852 2139 4160 2148
rect 4356 1442 4384 2790
rect 4540 2378 4568 3334
rect 5092 3126 5120 4422
rect 5184 3194 5212 5714
rect 5276 5370 5304 6190
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 5914 5580 6054
rect 6182 6012 6490 6021
rect 6182 6010 6188 6012
rect 6244 6010 6268 6012
rect 6324 6010 6348 6012
rect 6404 6010 6428 6012
rect 6484 6010 6490 6012
rect 6244 5958 6246 6010
rect 6426 5958 6428 6010
rect 6182 5956 6188 5958
rect 6244 5956 6268 5958
rect 6324 5956 6348 5958
rect 6404 5956 6428 5958
rect 6484 5956 6490 5958
rect 6182 5947 6490 5956
rect 6564 5914 6592 6802
rect 6842 6556 7150 6565
rect 6842 6554 6848 6556
rect 6904 6554 6928 6556
rect 6984 6554 7008 6556
rect 7064 6554 7088 6556
rect 7144 6554 7150 6556
rect 6904 6502 6906 6554
rect 7086 6502 7088 6554
rect 6842 6500 6848 6502
rect 6904 6500 6928 6502
rect 6984 6500 7008 6502
rect 7064 6500 7088 6502
rect 7144 6500 7150 6502
rect 6842 6491 7150 6500
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5347 5468 5655 5477
rect 5347 5466 5353 5468
rect 5409 5466 5433 5468
rect 5489 5466 5513 5468
rect 5569 5466 5593 5468
rect 5649 5466 5655 5468
rect 5409 5414 5411 5466
rect 5591 5414 5593 5466
rect 5347 5412 5353 5414
rect 5409 5412 5433 5414
rect 5489 5412 5513 5414
rect 5569 5412 5593 5414
rect 5649 5412 5655 5414
rect 5347 5403 5655 5412
rect 6104 5370 6132 5578
rect 7286 5536 7342 5545
rect 6842 5468 7150 5477
rect 7286 5471 7342 5480
rect 6842 5466 6848 5468
rect 6904 5466 6928 5468
rect 6984 5466 7008 5468
rect 7064 5466 7088 5468
rect 7144 5466 7150 5468
rect 6904 5414 6906 5466
rect 7086 5414 7088 5466
rect 6842 5412 6848 5414
rect 6904 5412 6928 5414
rect 6984 5412 7008 5414
rect 7064 5412 7088 5414
rect 7144 5412 7150 5414
rect 6842 5403 7150 5412
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 3738 5304 4422
rect 5347 4380 5655 4389
rect 5347 4378 5353 4380
rect 5409 4378 5433 4380
rect 5489 4378 5513 4380
rect 5569 4378 5593 4380
rect 5649 4378 5655 4380
rect 5409 4326 5411 4378
rect 5591 4326 5593 4378
rect 5347 4324 5353 4326
rect 5409 4324 5433 4326
rect 5489 4324 5513 4326
rect 5569 4324 5593 4326
rect 5649 4324 5655 4326
rect 5347 4315 5655 4324
rect 5736 4282 5764 5034
rect 5828 4758 5856 5034
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5920 4570 5948 5034
rect 5828 4542 5948 4570
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5828 4078 5856 4542
rect 6012 4486 6040 5102
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6104 4690 6132 4966
rect 6182 4924 6490 4933
rect 6182 4922 6188 4924
rect 6244 4922 6268 4924
rect 6324 4922 6348 4924
rect 6404 4922 6428 4924
rect 6484 4922 6490 4924
rect 6244 4870 6246 4922
rect 6426 4870 6428 4922
rect 6182 4868 6188 4870
rect 6244 4868 6268 4870
rect 6324 4868 6348 4870
rect 6404 4868 6428 4870
rect 6484 4868 6490 4870
rect 6182 4859 6490 4868
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5828 3466 5856 4014
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5347 3292 5655 3301
rect 5347 3290 5353 3292
rect 5409 3290 5433 3292
rect 5489 3290 5513 3292
rect 5569 3290 5593 3292
rect 5649 3290 5655 3292
rect 5409 3238 5411 3290
rect 5591 3238 5593 3290
rect 5347 3236 5353 3238
rect 5409 3236 5433 3238
rect 5489 3236 5513 3238
rect 5569 3236 5593 3238
rect 5649 3236 5655 3238
rect 5347 3227 5655 3236
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4687 2748 4995 2757
rect 4687 2746 4693 2748
rect 4749 2746 4773 2748
rect 4829 2746 4853 2748
rect 4909 2746 4933 2748
rect 4989 2746 4995 2748
rect 4749 2694 4751 2746
rect 4931 2694 4933 2746
rect 4687 2692 4693 2694
rect 4749 2692 4773 2694
rect 4829 2692 4853 2694
rect 4909 2692 4933 2694
rect 4989 2692 4995 2694
rect 4687 2683 4995 2692
rect 5184 2514 5212 3130
rect 5736 2514 5764 3334
rect 5828 2922 5856 3402
rect 6012 2990 6040 4422
rect 6842 4380 7150 4389
rect 6842 4378 6848 4380
rect 6904 4378 6928 4380
rect 6984 4378 7008 4380
rect 7064 4378 7088 4380
rect 7144 4378 7150 4380
rect 6904 4326 6906 4378
rect 7086 4326 7088 4378
rect 6842 4324 6848 4326
rect 6904 4324 6928 4326
rect 6984 4324 7008 4326
rect 7064 4324 7088 4326
rect 7144 4324 7150 4326
rect 6842 4315 7150 4324
rect 7300 4078 7328 5471
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 6182 3836 6490 3845
rect 6182 3834 6188 3836
rect 6244 3834 6268 3836
rect 6324 3834 6348 3836
rect 6404 3834 6428 3836
rect 6484 3834 6490 3836
rect 6244 3782 6246 3834
rect 6426 3782 6428 3834
rect 6182 3780 6188 3782
rect 6244 3780 6268 3782
rect 6324 3780 6348 3782
rect 6404 3780 6428 3782
rect 6484 3780 6490 3782
rect 6182 3771 6490 3780
rect 6842 3292 7150 3301
rect 6842 3290 6848 3292
rect 6904 3290 6928 3292
rect 6984 3290 7008 3292
rect 7064 3290 7088 3292
rect 7144 3290 7150 3292
rect 6904 3238 6906 3290
rect 7086 3238 7088 3290
rect 6842 3236 6848 3238
rect 6904 3236 6928 3238
rect 6984 3236 7008 3238
rect 7064 3236 7088 3238
rect 7144 3236 7150 3238
rect 6842 3227 7150 3236
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5828 2582 5856 2858
rect 6012 2650 6040 2926
rect 6182 2748 6490 2757
rect 6182 2746 6188 2748
rect 6244 2746 6268 2748
rect 6324 2746 6348 2748
rect 6404 2746 6428 2748
rect 6484 2746 6490 2748
rect 6244 2694 6246 2746
rect 6426 2694 6428 2746
rect 6182 2692 6188 2694
rect 6244 2692 6268 2694
rect 6324 2692 6348 2694
rect 6404 2692 6428 2694
rect 6484 2692 6490 2694
rect 6182 2683 6490 2692
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 5347 2204 5655 2213
rect 5347 2202 5353 2204
rect 5409 2202 5433 2204
rect 5489 2202 5513 2204
rect 5569 2202 5593 2204
rect 5649 2202 5655 2204
rect 5409 2150 5411 2202
rect 5591 2150 5593 2202
rect 5347 2148 5353 2150
rect 5409 2148 5433 2150
rect 5489 2148 5513 2150
rect 5569 2148 5593 2150
rect 5649 2148 5655 2150
rect 5347 2139 5655 2148
rect 6842 2204 7150 2213
rect 6842 2202 6848 2204
rect 6904 2202 6928 2204
rect 6984 2202 7008 2204
rect 7064 2202 7088 2204
rect 7144 2202 7150 2204
rect 6904 2150 6906 2202
rect 7086 2150 7088 2202
rect 6842 2148 6848 2150
rect 6904 2148 6928 2150
rect 6984 2148 7008 2150
rect 7064 2148 7088 2150
rect 7144 2148 7150 2150
rect 6842 2139 7150 2148
rect 4356 1414 4568 1442
rect 4540 800 4568 1414
rect 18 0 74 800
rect 4526 0 4582 800
rect 7208 785 7236 2314
rect 7194 776 7250 785
rect 7194 711 7250 720
<< via2 >>
rect 1398 9424 1454 9480
rect 1703 8186 1759 8188
rect 1783 8186 1839 8188
rect 1863 8186 1919 8188
rect 1943 8186 1999 8188
rect 1703 8134 1749 8186
rect 1749 8134 1759 8186
rect 1783 8134 1813 8186
rect 1813 8134 1825 8186
rect 1825 8134 1839 8186
rect 1863 8134 1877 8186
rect 1877 8134 1889 8186
rect 1889 8134 1919 8186
rect 1943 8134 1953 8186
rect 1953 8134 1999 8186
rect 1703 8132 1759 8134
rect 1783 8132 1839 8134
rect 1863 8132 1919 8134
rect 1943 8132 1999 8134
rect 3198 8186 3254 8188
rect 3278 8186 3334 8188
rect 3358 8186 3414 8188
rect 3438 8186 3494 8188
rect 3198 8134 3244 8186
rect 3244 8134 3254 8186
rect 3278 8134 3308 8186
rect 3308 8134 3320 8186
rect 3320 8134 3334 8186
rect 3358 8134 3372 8186
rect 3372 8134 3384 8186
rect 3384 8134 3414 8186
rect 3438 8134 3448 8186
rect 3448 8134 3494 8186
rect 3198 8132 3254 8134
rect 3278 8132 3334 8134
rect 3358 8132 3414 8134
rect 3438 8132 3494 8134
rect 4693 8186 4749 8188
rect 4773 8186 4829 8188
rect 4853 8186 4909 8188
rect 4933 8186 4989 8188
rect 4693 8134 4739 8186
rect 4739 8134 4749 8186
rect 4773 8134 4803 8186
rect 4803 8134 4815 8186
rect 4815 8134 4829 8186
rect 4853 8134 4867 8186
rect 4867 8134 4879 8186
rect 4879 8134 4909 8186
rect 4933 8134 4943 8186
rect 4943 8134 4989 8186
rect 4693 8132 4749 8134
rect 4773 8132 4829 8134
rect 4853 8132 4909 8134
rect 4933 8132 4989 8134
rect 6188 8186 6244 8188
rect 6268 8186 6324 8188
rect 6348 8186 6404 8188
rect 6428 8186 6484 8188
rect 6188 8134 6234 8186
rect 6234 8134 6244 8186
rect 6268 8134 6298 8186
rect 6298 8134 6310 8186
rect 6310 8134 6324 8186
rect 6348 8134 6362 8186
rect 6362 8134 6374 8186
rect 6374 8134 6404 8186
rect 6428 8134 6438 8186
rect 6438 8134 6484 8186
rect 6188 8132 6244 8134
rect 6268 8132 6324 8134
rect 6348 8132 6404 8134
rect 6428 8132 6484 8134
rect 1703 7098 1759 7100
rect 1783 7098 1839 7100
rect 1863 7098 1919 7100
rect 1943 7098 1999 7100
rect 1703 7046 1749 7098
rect 1749 7046 1759 7098
rect 1783 7046 1813 7098
rect 1813 7046 1825 7098
rect 1825 7046 1839 7098
rect 1863 7046 1877 7098
rect 1877 7046 1889 7098
rect 1889 7046 1919 7098
rect 1943 7046 1953 7098
rect 1953 7046 1999 7098
rect 1703 7044 1759 7046
rect 1783 7044 1839 7046
rect 1863 7044 1919 7046
rect 1943 7044 1999 7046
rect 1703 6010 1759 6012
rect 1783 6010 1839 6012
rect 1863 6010 1919 6012
rect 1943 6010 1999 6012
rect 1703 5958 1749 6010
rect 1749 5958 1759 6010
rect 1783 5958 1813 6010
rect 1813 5958 1825 6010
rect 1825 5958 1839 6010
rect 1863 5958 1877 6010
rect 1877 5958 1889 6010
rect 1889 5958 1919 6010
rect 1943 5958 1953 6010
rect 1953 5958 1999 6010
rect 1703 5956 1759 5958
rect 1783 5956 1839 5958
rect 1863 5956 1919 5958
rect 1943 5956 1999 5958
rect 2363 7642 2419 7644
rect 2443 7642 2499 7644
rect 2523 7642 2579 7644
rect 2603 7642 2659 7644
rect 2363 7590 2409 7642
rect 2409 7590 2419 7642
rect 2443 7590 2473 7642
rect 2473 7590 2485 7642
rect 2485 7590 2499 7642
rect 2523 7590 2537 7642
rect 2537 7590 2549 7642
rect 2549 7590 2579 7642
rect 2603 7590 2613 7642
rect 2613 7590 2659 7642
rect 2363 7588 2419 7590
rect 2443 7588 2499 7590
rect 2523 7588 2579 7590
rect 2603 7588 2659 7590
rect 2363 6554 2419 6556
rect 2443 6554 2499 6556
rect 2523 6554 2579 6556
rect 2603 6554 2659 6556
rect 2363 6502 2409 6554
rect 2409 6502 2419 6554
rect 2443 6502 2473 6554
rect 2473 6502 2485 6554
rect 2485 6502 2499 6554
rect 2523 6502 2537 6554
rect 2537 6502 2549 6554
rect 2549 6502 2579 6554
rect 2603 6502 2613 6554
rect 2613 6502 2659 6554
rect 2363 6500 2419 6502
rect 2443 6500 2499 6502
rect 2523 6500 2579 6502
rect 2603 6500 2659 6502
rect 3858 7642 3914 7644
rect 3938 7642 3994 7644
rect 4018 7642 4074 7644
rect 4098 7642 4154 7644
rect 3858 7590 3904 7642
rect 3904 7590 3914 7642
rect 3938 7590 3968 7642
rect 3968 7590 3980 7642
rect 3980 7590 3994 7642
rect 4018 7590 4032 7642
rect 4032 7590 4044 7642
rect 4044 7590 4074 7642
rect 4098 7590 4108 7642
rect 4108 7590 4154 7642
rect 3858 7588 3914 7590
rect 3938 7588 3994 7590
rect 4018 7588 4074 7590
rect 4098 7588 4154 7590
rect 5353 7642 5409 7644
rect 5433 7642 5489 7644
rect 5513 7642 5569 7644
rect 5593 7642 5649 7644
rect 5353 7590 5399 7642
rect 5399 7590 5409 7642
rect 5433 7590 5463 7642
rect 5463 7590 5475 7642
rect 5475 7590 5489 7642
rect 5513 7590 5527 7642
rect 5527 7590 5539 7642
rect 5539 7590 5569 7642
rect 5593 7590 5603 7642
rect 5603 7590 5649 7642
rect 5353 7588 5409 7590
rect 5433 7588 5489 7590
rect 5513 7588 5569 7590
rect 5593 7588 5649 7590
rect 3198 7098 3254 7100
rect 3278 7098 3334 7100
rect 3358 7098 3414 7100
rect 3438 7098 3494 7100
rect 3198 7046 3244 7098
rect 3244 7046 3254 7098
rect 3278 7046 3308 7098
rect 3308 7046 3320 7098
rect 3320 7046 3334 7098
rect 3358 7046 3372 7098
rect 3372 7046 3384 7098
rect 3384 7046 3414 7098
rect 3438 7046 3448 7098
rect 3448 7046 3494 7098
rect 3198 7044 3254 7046
rect 3278 7044 3334 7046
rect 3358 7044 3414 7046
rect 3438 7044 3494 7046
rect 4693 7098 4749 7100
rect 4773 7098 4829 7100
rect 4853 7098 4909 7100
rect 4933 7098 4989 7100
rect 4693 7046 4739 7098
rect 4739 7046 4749 7098
rect 4773 7046 4803 7098
rect 4803 7046 4815 7098
rect 4815 7046 4829 7098
rect 4853 7046 4867 7098
rect 4867 7046 4879 7098
rect 4879 7046 4909 7098
rect 4933 7046 4943 7098
rect 4943 7046 4989 7098
rect 4693 7044 4749 7046
rect 4773 7044 4829 7046
rect 4853 7044 4909 7046
rect 4933 7044 4989 7046
rect 6848 7642 6904 7644
rect 6928 7642 6984 7644
rect 7008 7642 7064 7644
rect 7088 7642 7144 7644
rect 6848 7590 6894 7642
rect 6894 7590 6904 7642
rect 6928 7590 6958 7642
rect 6958 7590 6970 7642
rect 6970 7590 6984 7642
rect 7008 7590 7022 7642
rect 7022 7590 7034 7642
rect 7034 7590 7064 7642
rect 7088 7590 7098 7642
rect 7098 7590 7144 7642
rect 6848 7588 6904 7590
rect 6928 7588 6984 7590
rect 7008 7588 7064 7590
rect 7088 7588 7144 7590
rect 6188 7098 6244 7100
rect 6268 7098 6324 7100
rect 6348 7098 6404 7100
rect 6428 7098 6484 7100
rect 6188 7046 6234 7098
rect 6234 7046 6244 7098
rect 6268 7046 6298 7098
rect 6298 7046 6310 7098
rect 6310 7046 6324 7098
rect 6348 7046 6362 7098
rect 6362 7046 6374 7098
rect 6374 7046 6404 7098
rect 6428 7046 6438 7098
rect 6438 7046 6484 7098
rect 6188 7044 6244 7046
rect 6268 7044 6324 7046
rect 6348 7044 6404 7046
rect 6428 7044 6484 7046
rect 3858 6554 3914 6556
rect 3938 6554 3994 6556
rect 4018 6554 4074 6556
rect 4098 6554 4154 6556
rect 3858 6502 3904 6554
rect 3904 6502 3914 6554
rect 3938 6502 3968 6554
rect 3968 6502 3980 6554
rect 3980 6502 3994 6554
rect 4018 6502 4032 6554
rect 4032 6502 4044 6554
rect 4044 6502 4074 6554
rect 4098 6502 4108 6554
rect 4108 6502 4154 6554
rect 3858 6500 3914 6502
rect 3938 6500 3994 6502
rect 4018 6500 4074 6502
rect 4098 6500 4154 6502
rect 3198 6010 3254 6012
rect 3278 6010 3334 6012
rect 3358 6010 3414 6012
rect 3438 6010 3494 6012
rect 3198 5958 3244 6010
rect 3244 5958 3254 6010
rect 3278 5958 3308 6010
rect 3308 5958 3320 6010
rect 3320 5958 3334 6010
rect 3358 5958 3372 6010
rect 3372 5958 3384 6010
rect 3384 5958 3414 6010
rect 3438 5958 3448 6010
rect 3448 5958 3494 6010
rect 3198 5956 3254 5958
rect 3278 5956 3334 5958
rect 3358 5956 3414 5958
rect 3438 5956 3494 5958
rect 4693 6010 4749 6012
rect 4773 6010 4829 6012
rect 4853 6010 4909 6012
rect 4933 6010 4989 6012
rect 4693 5958 4739 6010
rect 4739 5958 4749 6010
rect 4773 5958 4803 6010
rect 4803 5958 4815 6010
rect 4815 5958 4829 6010
rect 4853 5958 4867 6010
rect 4867 5958 4879 6010
rect 4879 5958 4909 6010
rect 4933 5958 4943 6010
rect 4943 5958 4989 6010
rect 4693 5956 4749 5958
rect 4773 5956 4829 5958
rect 4853 5956 4909 5958
rect 4933 5956 4989 5958
rect 1703 4922 1759 4924
rect 1783 4922 1839 4924
rect 1863 4922 1919 4924
rect 1943 4922 1999 4924
rect 1703 4870 1749 4922
rect 1749 4870 1759 4922
rect 1783 4870 1813 4922
rect 1813 4870 1825 4922
rect 1825 4870 1839 4922
rect 1863 4870 1877 4922
rect 1877 4870 1889 4922
rect 1889 4870 1919 4922
rect 1943 4870 1953 4922
rect 1953 4870 1999 4922
rect 1703 4868 1759 4870
rect 1783 4868 1839 4870
rect 1863 4868 1919 4870
rect 1943 4868 1999 4870
rect 938 4800 994 4856
rect 1703 3834 1759 3836
rect 1783 3834 1839 3836
rect 1863 3834 1919 3836
rect 1943 3834 1999 3836
rect 1703 3782 1749 3834
rect 1749 3782 1759 3834
rect 1783 3782 1813 3834
rect 1813 3782 1825 3834
rect 1825 3782 1839 3834
rect 1863 3782 1877 3834
rect 1877 3782 1889 3834
rect 1889 3782 1919 3834
rect 1943 3782 1953 3834
rect 1953 3782 1999 3834
rect 1703 3780 1759 3782
rect 1783 3780 1839 3782
rect 1863 3780 1919 3782
rect 1943 3780 1999 3782
rect 2363 5466 2419 5468
rect 2443 5466 2499 5468
rect 2523 5466 2579 5468
rect 2603 5466 2659 5468
rect 2363 5414 2409 5466
rect 2409 5414 2419 5466
rect 2443 5414 2473 5466
rect 2473 5414 2485 5466
rect 2485 5414 2499 5466
rect 2523 5414 2537 5466
rect 2537 5414 2549 5466
rect 2549 5414 2579 5466
rect 2603 5414 2613 5466
rect 2613 5414 2659 5466
rect 2363 5412 2419 5414
rect 2443 5412 2499 5414
rect 2523 5412 2579 5414
rect 2603 5412 2659 5414
rect 2363 4378 2419 4380
rect 2443 4378 2499 4380
rect 2523 4378 2579 4380
rect 2603 4378 2659 4380
rect 2363 4326 2409 4378
rect 2409 4326 2419 4378
rect 2443 4326 2473 4378
rect 2473 4326 2485 4378
rect 2485 4326 2499 4378
rect 2523 4326 2537 4378
rect 2537 4326 2549 4378
rect 2549 4326 2579 4378
rect 2603 4326 2613 4378
rect 2613 4326 2659 4378
rect 2363 4324 2419 4326
rect 2443 4324 2499 4326
rect 2523 4324 2579 4326
rect 2603 4324 2659 4326
rect 2363 3290 2419 3292
rect 2443 3290 2499 3292
rect 2523 3290 2579 3292
rect 2603 3290 2659 3292
rect 2363 3238 2409 3290
rect 2409 3238 2419 3290
rect 2443 3238 2473 3290
rect 2473 3238 2485 3290
rect 2485 3238 2499 3290
rect 2523 3238 2537 3290
rect 2537 3238 2549 3290
rect 2549 3238 2579 3290
rect 2603 3238 2613 3290
rect 2613 3238 2659 3290
rect 2363 3236 2419 3238
rect 2443 3236 2499 3238
rect 2523 3236 2579 3238
rect 2603 3236 2659 3238
rect 3858 5466 3914 5468
rect 3938 5466 3994 5468
rect 4018 5466 4074 5468
rect 4098 5466 4154 5468
rect 3858 5414 3904 5466
rect 3904 5414 3914 5466
rect 3938 5414 3968 5466
rect 3968 5414 3980 5466
rect 3980 5414 3994 5466
rect 4018 5414 4032 5466
rect 4032 5414 4044 5466
rect 4044 5414 4074 5466
rect 4098 5414 4108 5466
rect 4108 5414 4154 5466
rect 3858 5412 3914 5414
rect 3938 5412 3994 5414
rect 4018 5412 4074 5414
rect 4098 5412 4154 5414
rect 3198 4922 3254 4924
rect 3278 4922 3334 4924
rect 3358 4922 3414 4924
rect 3438 4922 3494 4924
rect 3198 4870 3244 4922
rect 3244 4870 3254 4922
rect 3278 4870 3308 4922
rect 3308 4870 3320 4922
rect 3320 4870 3334 4922
rect 3358 4870 3372 4922
rect 3372 4870 3384 4922
rect 3384 4870 3414 4922
rect 3438 4870 3448 4922
rect 3448 4870 3494 4922
rect 3198 4868 3254 4870
rect 3278 4868 3334 4870
rect 3358 4868 3414 4870
rect 3438 4868 3494 4870
rect 5353 6554 5409 6556
rect 5433 6554 5489 6556
rect 5513 6554 5569 6556
rect 5593 6554 5649 6556
rect 5353 6502 5399 6554
rect 5399 6502 5409 6554
rect 5433 6502 5463 6554
rect 5463 6502 5475 6554
rect 5475 6502 5489 6554
rect 5513 6502 5527 6554
rect 5527 6502 5539 6554
rect 5539 6502 5569 6554
rect 5593 6502 5603 6554
rect 5603 6502 5649 6554
rect 5353 6500 5409 6502
rect 5433 6500 5489 6502
rect 5513 6500 5569 6502
rect 5593 6500 5649 6502
rect 4693 4922 4749 4924
rect 4773 4922 4829 4924
rect 4853 4922 4909 4924
rect 4933 4922 4989 4924
rect 4693 4870 4739 4922
rect 4739 4870 4749 4922
rect 4773 4870 4803 4922
rect 4803 4870 4815 4922
rect 4815 4870 4829 4922
rect 4853 4870 4867 4922
rect 4867 4870 4879 4922
rect 4879 4870 4909 4922
rect 4933 4870 4943 4922
rect 4943 4870 4989 4922
rect 4693 4868 4749 4870
rect 4773 4868 4829 4870
rect 4853 4868 4909 4870
rect 4933 4868 4989 4870
rect 3858 4378 3914 4380
rect 3938 4378 3994 4380
rect 4018 4378 4074 4380
rect 4098 4378 4154 4380
rect 3858 4326 3904 4378
rect 3904 4326 3914 4378
rect 3938 4326 3968 4378
rect 3968 4326 3980 4378
rect 3980 4326 3994 4378
rect 4018 4326 4032 4378
rect 4032 4326 4044 4378
rect 4044 4326 4074 4378
rect 4098 4326 4108 4378
rect 4108 4326 4154 4378
rect 3858 4324 3914 4326
rect 3938 4324 3994 4326
rect 4018 4324 4074 4326
rect 4098 4324 4154 4326
rect 3198 3834 3254 3836
rect 3278 3834 3334 3836
rect 3358 3834 3414 3836
rect 3438 3834 3494 3836
rect 3198 3782 3244 3834
rect 3244 3782 3254 3834
rect 3278 3782 3308 3834
rect 3308 3782 3320 3834
rect 3320 3782 3334 3834
rect 3358 3782 3372 3834
rect 3372 3782 3384 3834
rect 3384 3782 3414 3834
rect 3438 3782 3448 3834
rect 3448 3782 3494 3834
rect 3198 3780 3254 3782
rect 3278 3780 3334 3782
rect 3358 3780 3414 3782
rect 3438 3780 3494 3782
rect 4693 3834 4749 3836
rect 4773 3834 4829 3836
rect 4853 3834 4909 3836
rect 4933 3834 4989 3836
rect 4693 3782 4739 3834
rect 4739 3782 4749 3834
rect 4773 3782 4803 3834
rect 4803 3782 4815 3834
rect 4815 3782 4829 3834
rect 4853 3782 4867 3834
rect 4867 3782 4879 3834
rect 4879 3782 4909 3834
rect 4933 3782 4943 3834
rect 4943 3782 4989 3834
rect 4693 3780 4749 3782
rect 4773 3780 4829 3782
rect 4853 3780 4909 3782
rect 4933 3780 4989 3782
rect 3858 3290 3914 3292
rect 3938 3290 3994 3292
rect 4018 3290 4074 3292
rect 4098 3290 4154 3292
rect 3858 3238 3904 3290
rect 3904 3238 3914 3290
rect 3938 3238 3968 3290
rect 3968 3238 3980 3290
rect 3980 3238 3994 3290
rect 4018 3238 4032 3290
rect 4032 3238 4044 3290
rect 4044 3238 4074 3290
rect 4098 3238 4108 3290
rect 4108 3238 4154 3290
rect 3858 3236 3914 3238
rect 3938 3236 3994 3238
rect 4018 3236 4074 3238
rect 4098 3236 4154 3238
rect 18 2896 74 2952
rect 2870 2896 2926 2952
rect 1703 2746 1759 2748
rect 1783 2746 1839 2748
rect 1863 2746 1919 2748
rect 1943 2746 1999 2748
rect 1703 2694 1749 2746
rect 1749 2694 1759 2746
rect 1783 2694 1813 2746
rect 1813 2694 1825 2746
rect 1825 2694 1839 2746
rect 1863 2694 1877 2746
rect 1877 2694 1889 2746
rect 1889 2694 1919 2746
rect 1943 2694 1953 2746
rect 1953 2694 1999 2746
rect 1703 2692 1759 2694
rect 1783 2692 1839 2694
rect 1863 2692 1919 2694
rect 1943 2692 1999 2694
rect 3198 2746 3254 2748
rect 3278 2746 3334 2748
rect 3358 2746 3414 2748
rect 3438 2746 3494 2748
rect 3198 2694 3244 2746
rect 3244 2694 3254 2746
rect 3278 2694 3308 2746
rect 3308 2694 3320 2746
rect 3320 2694 3334 2746
rect 3358 2694 3372 2746
rect 3372 2694 3384 2746
rect 3384 2694 3414 2746
rect 3438 2694 3448 2746
rect 3448 2694 3494 2746
rect 3198 2692 3254 2694
rect 3278 2692 3334 2694
rect 3358 2692 3414 2694
rect 3438 2692 3494 2694
rect 2363 2202 2419 2204
rect 2443 2202 2499 2204
rect 2523 2202 2579 2204
rect 2603 2202 2659 2204
rect 2363 2150 2409 2202
rect 2409 2150 2419 2202
rect 2443 2150 2473 2202
rect 2473 2150 2485 2202
rect 2485 2150 2499 2202
rect 2523 2150 2537 2202
rect 2537 2150 2549 2202
rect 2549 2150 2579 2202
rect 2603 2150 2613 2202
rect 2613 2150 2659 2202
rect 2363 2148 2419 2150
rect 2443 2148 2499 2150
rect 2523 2148 2579 2150
rect 2603 2148 2659 2150
rect 3858 2202 3914 2204
rect 3938 2202 3994 2204
rect 4018 2202 4074 2204
rect 4098 2202 4154 2204
rect 3858 2150 3904 2202
rect 3904 2150 3914 2202
rect 3938 2150 3968 2202
rect 3968 2150 3980 2202
rect 3980 2150 3994 2202
rect 4018 2150 4032 2202
rect 4032 2150 4044 2202
rect 4044 2150 4074 2202
rect 4098 2150 4108 2202
rect 4108 2150 4154 2202
rect 3858 2148 3914 2150
rect 3938 2148 3994 2150
rect 4018 2148 4074 2150
rect 4098 2148 4154 2150
rect 6188 6010 6244 6012
rect 6268 6010 6324 6012
rect 6348 6010 6404 6012
rect 6428 6010 6484 6012
rect 6188 5958 6234 6010
rect 6234 5958 6244 6010
rect 6268 5958 6298 6010
rect 6298 5958 6310 6010
rect 6310 5958 6324 6010
rect 6348 5958 6362 6010
rect 6362 5958 6374 6010
rect 6374 5958 6404 6010
rect 6428 5958 6438 6010
rect 6438 5958 6484 6010
rect 6188 5956 6244 5958
rect 6268 5956 6324 5958
rect 6348 5956 6404 5958
rect 6428 5956 6484 5958
rect 6848 6554 6904 6556
rect 6928 6554 6984 6556
rect 7008 6554 7064 6556
rect 7088 6554 7144 6556
rect 6848 6502 6894 6554
rect 6894 6502 6904 6554
rect 6928 6502 6958 6554
rect 6958 6502 6970 6554
rect 6970 6502 6984 6554
rect 7008 6502 7022 6554
rect 7022 6502 7034 6554
rect 7034 6502 7064 6554
rect 7088 6502 7098 6554
rect 7098 6502 7144 6554
rect 6848 6500 6904 6502
rect 6928 6500 6984 6502
rect 7008 6500 7064 6502
rect 7088 6500 7144 6502
rect 5353 5466 5409 5468
rect 5433 5466 5489 5468
rect 5513 5466 5569 5468
rect 5593 5466 5649 5468
rect 5353 5414 5399 5466
rect 5399 5414 5409 5466
rect 5433 5414 5463 5466
rect 5463 5414 5475 5466
rect 5475 5414 5489 5466
rect 5513 5414 5527 5466
rect 5527 5414 5539 5466
rect 5539 5414 5569 5466
rect 5593 5414 5603 5466
rect 5603 5414 5649 5466
rect 5353 5412 5409 5414
rect 5433 5412 5489 5414
rect 5513 5412 5569 5414
rect 5593 5412 5649 5414
rect 7286 5480 7342 5536
rect 6848 5466 6904 5468
rect 6928 5466 6984 5468
rect 7008 5466 7064 5468
rect 7088 5466 7144 5468
rect 6848 5414 6894 5466
rect 6894 5414 6904 5466
rect 6928 5414 6958 5466
rect 6958 5414 6970 5466
rect 6970 5414 6984 5466
rect 7008 5414 7022 5466
rect 7022 5414 7034 5466
rect 7034 5414 7064 5466
rect 7088 5414 7098 5466
rect 7098 5414 7144 5466
rect 6848 5412 6904 5414
rect 6928 5412 6984 5414
rect 7008 5412 7064 5414
rect 7088 5412 7144 5414
rect 5353 4378 5409 4380
rect 5433 4378 5489 4380
rect 5513 4378 5569 4380
rect 5593 4378 5649 4380
rect 5353 4326 5399 4378
rect 5399 4326 5409 4378
rect 5433 4326 5463 4378
rect 5463 4326 5475 4378
rect 5475 4326 5489 4378
rect 5513 4326 5527 4378
rect 5527 4326 5539 4378
rect 5539 4326 5569 4378
rect 5593 4326 5603 4378
rect 5603 4326 5649 4378
rect 5353 4324 5409 4326
rect 5433 4324 5489 4326
rect 5513 4324 5569 4326
rect 5593 4324 5649 4326
rect 6188 4922 6244 4924
rect 6268 4922 6324 4924
rect 6348 4922 6404 4924
rect 6428 4922 6484 4924
rect 6188 4870 6234 4922
rect 6234 4870 6244 4922
rect 6268 4870 6298 4922
rect 6298 4870 6310 4922
rect 6310 4870 6324 4922
rect 6348 4870 6362 4922
rect 6362 4870 6374 4922
rect 6374 4870 6404 4922
rect 6428 4870 6438 4922
rect 6438 4870 6484 4922
rect 6188 4868 6244 4870
rect 6268 4868 6324 4870
rect 6348 4868 6404 4870
rect 6428 4868 6484 4870
rect 5353 3290 5409 3292
rect 5433 3290 5489 3292
rect 5513 3290 5569 3292
rect 5593 3290 5649 3292
rect 5353 3238 5399 3290
rect 5399 3238 5409 3290
rect 5433 3238 5463 3290
rect 5463 3238 5475 3290
rect 5475 3238 5489 3290
rect 5513 3238 5527 3290
rect 5527 3238 5539 3290
rect 5539 3238 5569 3290
rect 5593 3238 5603 3290
rect 5603 3238 5649 3290
rect 5353 3236 5409 3238
rect 5433 3236 5489 3238
rect 5513 3236 5569 3238
rect 5593 3236 5649 3238
rect 4693 2746 4749 2748
rect 4773 2746 4829 2748
rect 4853 2746 4909 2748
rect 4933 2746 4989 2748
rect 4693 2694 4739 2746
rect 4739 2694 4749 2746
rect 4773 2694 4803 2746
rect 4803 2694 4815 2746
rect 4815 2694 4829 2746
rect 4853 2694 4867 2746
rect 4867 2694 4879 2746
rect 4879 2694 4909 2746
rect 4933 2694 4943 2746
rect 4943 2694 4989 2746
rect 4693 2692 4749 2694
rect 4773 2692 4829 2694
rect 4853 2692 4909 2694
rect 4933 2692 4989 2694
rect 6848 4378 6904 4380
rect 6928 4378 6984 4380
rect 7008 4378 7064 4380
rect 7088 4378 7144 4380
rect 6848 4326 6894 4378
rect 6894 4326 6904 4378
rect 6928 4326 6958 4378
rect 6958 4326 6970 4378
rect 6970 4326 6984 4378
rect 7008 4326 7022 4378
rect 7022 4326 7034 4378
rect 7034 4326 7064 4378
rect 7088 4326 7098 4378
rect 7098 4326 7144 4378
rect 6848 4324 6904 4326
rect 6928 4324 6984 4326
rect 7008 4324 7064 4326
rect 7088 4324 7144 4326
rect 6188 3834 6244 3836
rect 6268 3834 6324 3836
rect 6348 3834 6404 3836
rect 6428 3834 6484 3836
rect 6188 3782 6234 3834
rect 6234 3782 6244 3834
rect 6268 3782 6298 3834
rect 6298 3782 6310 3834
rect 6310 3782 6324 3834
rect 6348 3782 6362 3834
rect 6362 3782 6374 3834
rect 6374 3782 6404 3834
rect 6428 3782 6438 3834
rect 6438 3782 6484 3834
rect 6188 3780 6244 3782
rect 6268 3780 6324 3782
rect 6348 3780 6404 3782
rect 6428 3780 6484 3782
rect 6848 3290 6904 3292
rect 6928 3290 6984 3292
rect 7008 3290 7064 3292
rect 7088 3290 7144 3292
rect 6848 3238 6894 3290
rect 6894 3238 6904 3290
rect 6928 3238 6958 3290
rect 6958 3238 6970 3290
rect 6970 3238 6984 3290
rect 7008 3238 7022 3290
rect 7022 3238 7034 3290
rect 7034 3238 7064 3290
rect 7088 3238 7098 3290
rect 7098 3238 7144 3290
rect 6848 3236 6904 3238
rect 6928 3236 6984 3238
rect 7008 3236 7064 3238
rect 7088 3236 7144 3238
rect 6188 2746 6244 2748
rect 6268 2746 6324 2748
rect 6348 2746 6404 2748
rect 6428 2746 6484 2748
rect 6188 2694 6234 2746
rect 6234 2694 6244 2746
rect 6268 2694 6298 2746
rect 6298 2694 6310 2746
rect 6310 2694 6324 2746
rect 6348 2694 6362 2746
rect 6362 2694 6374 2746
rect 6374 2694 6404 2746
rect 6428 2694 6438 2746
rect 6438 2694 6484 2746
rect 6188 2692 6244 2694
rect 6268 2692 6324 2694
rect 6348 2692 6404 2694
rect 6428 2692 6484 2694
rect 5353 2202 5409 2204
rect 5433 2202 5489 2204
rect 5513 2202 5569 2204
rect 5593 2202 5649 2204
rect 5353 2150 5399 2202
rect 5399 2150 5409 2202
rect 5433 2150 5463 2202
rect 5463 2150 5475 2202
rect 5475 2150 5489 2202
rect 5513 2150 5527 2202
rect 5527 2150 5539 2202
rect 5539 2150 5569 2202
rect 5593 2150 5603 2202
rect 5603 2150 5649 2202
rect 5353 2148 5409 2150
rect 5433 2148 5489 2150
rect 5513 2148 5569 2150
rect 5593 2148 5649 2150
rect 6848 2202 6904 2204
rect 6928 2202 6984 2204
rect 7008 2202 7064 2204
rect 7088 2202 7144 2204
rect 6848 2150 6894 2202
rect 6894 2150 6904 2202
rect 6928 2150 6958 2202
rect 6958 2150 6970 2202
rect 6970 2150 6984 2202
rect 7008 2150 7022 2202
rect 7022 2150 7034 2202
rect 7034 2150 7064 2202
rect 7088 2150 7098 2202
rect 7098 2150 7144 2202
rect 6848 2148 6904 2150
rect 6928 2148 6984 2150
rect 7008 2148 7064 2150
rect 7088 2148 7144 2150
rect 7194 720 7250 776
<< metal3 >>
rect 0 9618 800 9648
rect 0 9558 1042 9618
rect 0 9528 800 9558
rect 982 9482 1042 9558
rect 1393 9482 1459 9485
rect 982 9480 1459 9482
rect 982 9424 1398 9480
rect 1454 9424 1459 9480
rect 982 9422 1459 9424
rect 1393 9419 1459 9422
rect 1693 8192 2009 8193
rect 1693 8128 1699 8192
rect 1763 8128 1779 8192
rect 1843 8128 1859 8192
rect 1923 8128 1939 8192
rect 2003 8128 2009 8192
rect 1693 8127 2009 8128
rect 3188 8192 3504 8193
rect 3188 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3434 8192
rect 3498 8128 3504 8192
rect 3188 8127 3504 8128
rect 4683 8192 4999 8193
rect 4683 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4929 8192
rect 4993 8128 4999 8192
rect 4683 8127 4999 8128
rect 6178 8192 6494 8193
rect 6178 8128 6184 8192
rect 6248 8128 6264 8192
rect 6328 8128 6344 8192
rect 6408 8128 6424 8192
rect 6488 8128 6494 8192
rect 6178 8127 6494 8128
rect 2353 7648 2669 7649
rect 2353 7584 2359 7648
rect 2423 7584 2439 7648
rect 2503 7584 2519 7648
rect 2583 7584 2599 7648
rect 2663 7584 2669 7648
rect 2353 7583 2669 7584
rect 3848 7648 4164 7649
rect 3848 7584 3854 7648
rect 3918 7584 3934 7648
rect 3998 7584 4014 7648
rect 4078 7584 4094 7648
rect 4158 7584 4164 7648
rect 3848 7583 4164 7584
rect 5343 7648 5659 7649
rect 5343 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5589 7648
rect 5653 7584 5659 7648
rect 5343 7583 5659 7584
rect 6838 7648 7154 7649
rect 6838 7584 6844 7648
rect 6908 7584 6924 7648
rect 6988 7584 7004 7648
rect 7068 7584 7084 7648
rect 7148 7584 7154 7648
rect 6838 7583 7154 7584
rect 1693 7104 2009 7105
rect 1693 7040 1699 7104
rect 1763 7040 1779 7104
rect 1843 7040 1859 7104
rect 1923 7040 1939 7104
rect 2003 7040 2009 7104
rect 1693 7039 2009 7040
rect 3188 7104 3504 7105
rect 3188 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3434 7104
rect 3498 7040 3504 7104
rect 3188 7039 3504 7040
rect 4683 7104 4999 7105
rect 4683 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4929 7104
rect 4993 7040 4999 7104
rect 4683 7039 4999 7040
rect 6178 7104 6494 7105
rect 6178 7040 6184 7104
rect 6248 7040 6264 7104
rect 6328 7040 6344 7104
rect 6408 7040 6424 7104
rect 6488 7040 6494 7104
rect 6178 7039 6494 7040
rect 2353 6560 2669 6561
rect 2353 6496 2359 6560
rect 2423 6496 2439 6560
rect 2503 6496 2519 6560
rect 2583 6496 2599 6560
rect 2663 6496 2669 6560
rect 2353 6495 2669 6496
rect 3848 6560 4164 6561
rect 3848 6496 3854 6560
rect 3918 6496 3934 6560
rect 3998 6496 4014 6560
rect 4078 6496 4094 6560
rect 4158 6496 4164 6560
rect 3848 6495 4164 6496
rect 5343 6560 5659 6561
rect 5343 6496 5349 6560
rect 5413 6496 5429 6560
rect 5493 6496 5509 6560
rect 5573 6496 5589 6560
rect 5653 6496 5659 6560
rect 5343 6495 5659 6496
rect 6838 6560 7154 6561
rect 6838 6496 6844 6560
rect 6908 6496 6924 6560
rect 6988 6496 7004 6560
rect 7068 6496 7084 6560
rect 7148 6496 7154 6560
rect 6838 6495 7154 6496
rect 1693 6016 2009 6017
rect 1693 5952 1699 6016
rect 1763 5952 1779 6016
rect 1843 5952 1859 6016
rect 1923 5952 1939 6016
rect 2003 5952 2009 6016
rect 1693 5951 2009 5952
rect 3188 6016 3504 6017
rect 3188 5952 3194 6016
rect 3258 5952 3274 6016
rect 3338 5952 3354 6016
rect 3418 5952 3434 6016
rect 3498 5952 3504 6016
rect 3188 5951 3504 5952
rect 4683 6016 4999 6017
rect 4683 5952 4689 6016
rect 4753 5952 4769 6016
rect 4833 5952 4849 6016
rect 4913 5952 4929 6016
rect 4993 5952 4999 6016
rect 4683 5951 4999 5952
rect 6178 6016 6494 6017
rect 6178 5952 6184 6016
rect 6248 5952 6264 6016
rect 6328 5952 6344 6016
rect 6408 5952 6424 6016
rect 6488 5952 6494 6016
rect 6178 5951 6494 5952
rect 7281 5538 7347 5541
rect 7411 5538 8211 5568
rect 7281 5536 8211 5538
rect 7281 5480 7286 5536
rect 7342 5480 8211 5536
rect 7281 5478 8211 5480
rect 7281 5475 7347 5478
rect 2353 5472 2669 5473
rect 2353 5408 2359 5472
rect 2423 5408 2439 5472
rect 2503 5408 2519 5472
rect 2583 5408 2599 5472
rect 2663 5408 2669 5472
rect 2353 5407 2669 5408
rect 3848 5472 4164 5473
rect 3848 5408 3854 5472
rect 3918 5408 3934 5472
rect 3998 5408 4014 5472
rect 4078 5408 4094 5472
rect 4158 5408 4164 5472
rect 3848 5407 4164 5408
rect 5343 5472 5659 5473
rect 5343 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5589 5472
rect 5653 5408 5659 5472
rect 5343 5407 5659 5408
rect 6838 5472 7154 5473
rect 6838 5408 6844 5472
rect 6908 5408 6924 5472
rect 6988 5408 7004 5472
rect 7068 5408 7084 5472
rect 7148 5408 7154 5472
rect 7411 5448 8211 5478
rect 6838 5407 7154 5408
rect 1693 4928 2009 4929
rect 0 4858 800 4888
rect 1693 4864 1699 4928
rect 1763 4864 1779 4928
rect 1843 4864 1859 4928
rect 1923 4864 1939 4928
rect 2003 4864 2009 4928
rect 1693 4863 2009 4864
rect 3188 4928 3504 4929
rect 3188 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3434 4928
rect 3498 4864 3504 4928
rect 3188 4863 3504 4864
rect 4683 4928 4999 4929
rect 4683 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4929 4928
rect 4993 4864 4999 4928
rect 4683 4863 4999 4864
rect 6178 4928 6494 4929
rect 6178 4864 6184 4928
rect 6248 4864 6264 4928
rect 6328 4864 6344 4928
rect 6408 4864 6424 4928
rect 6488 4864 6494 4928
rect 6178 4863 6494 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 2353 4384 2669 4385
rect 2353 4320 2359 4384
rect 2423 4320 2439 4384
rect 2503 4320 2519 4384
rect 2583 4320 2599 4384
rect 2663 4320 2669 4384
rect 2353 4319 2669 4320
rect 3848 4384 4164 4385
rect 3848 4320 3854 4384
rect 3918 4320 3934 4384
rect 3998 4320 4014 4384
rect 4078 4320 4094 4384
rect 4158 4320 4164 4384
rect 3848 4319 4164 4320
rect 5343 4384 5659 4385
rect 5343 4320 5349 4384
rect 5413 4320 5429 4384
rect 5493 4320 5509 4384
rect 5573 4320 5589 4384
rect 5653 4320 5659 4384
rect 5343 4319 5659 4320
rect 6838 4384 7154 4385
rect 6838 4320 6844 4384
rect 6908 4320 6924 4384
rect 6988 4320 7004 4384
rect 7068 4320 7084 4384
rect 7148 4320 7154 4384
rect 6838 4319 7154 4320
rect 1693 3840 2009 3841
rect 1693 3776 1699 3840
rect 1763 3776 1779 3840
rect 1843 3776 1859 3840
rect 1923 3776 1939 3840
rect 2003 3776 2009 3840
rect 1693 3775 2009 3776
rect 3188 3840 3504 3841
rect 3188 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3434 3840
rect 3498 3776 3504 3840
rect 3188 3775 3504 3776
rect 4683 3840 4999 3841
rect 4683 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4929 3840
rect 4993 3776 4999 3840
rect 4683 3775 4999 3776
rect 6178 3840 6494 3841
rect 6178 3776 6184 3840
rect 6248 3776 6264 3840
rect 6328 3776 6344 3840
rect 6408 3776 6424 3840
rect 6488 3776 6494 3840
rect 6178 3775 6494 3776
rect 2353 3296 2669 3297
rect 2353 3232 2359 3296
rect 2423 3232 2439 3296
rect 2503 3232 2519 3296
rect 2583 3232 2599 3296
rect 2663 3232 2669 3296
rect 2353 3231 2669 3232
rect 3848 3296 4164 3297
rect 3848 3232 3854 3296
rect 3918 3232 3934 3296
rect 3998 3232 4014 3296
rect 4078 3232 4094 3296
rect 4158 3232 4164 3296
rect 3848 3231 4164 3232
rect 5343 3296 5659 3297
rect 5343 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5589 3296
rect 5653 3232 5659 3296
rect 5343 3231 5659 3232
rect 6838 3296 7154 3297
rect 6838 3232 6844 3296
rect 6908 3232 6924 3296
rect 6988 3232 7004 3296
rect 7068 3232 7084 3296
rect 7148 3232 7154 3296
rect 6838 3231 7154 3232
rect 13 2954 79 2957
rect 2865 2954 2931 2957
rect 13 2952 2931 2954
rect 13 2896 18 2952
rect 74 2896 2870 2952
rect 2926 2896 2931 2952
rect 13 2894 2931 2896
rect 13 2891 79 2894
rect 2865 2891 2931 2894
rect 1693 2752 2009 2753
rect 1693 2688 1699 2752
rect 1763 2688 1779 2752
rect 1843 2688 1859 2752
rect 1923 2688 1939 2752
rect 2003 2688 2009 2752
rect 1693 2687 2009 2688
rect 3188 2752 3504 2753
rect 3188 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3434 2752
rect 3498 2688 3504 2752
rect 3188 2687 3504 2688
rect 4683 2752 4999 2753
rect 4683 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4929 2752
rect 4993 2688 4999 2752
rect 4683 2687 4999 2688
rect 6178 2752 6494 2753
rect 6178 2688 6184 2752
rect 6248 2688 6264 2752
rect 6328 2688 6344 2752
rect 6408 2688 6424 2752
rect 6488 2688 6494 2752
rect 6178 2687 6494 2688
rect 2353 2208 2669 2209
rect 2353 2144 2359 2208
rect 2423 2144 2439 2208
rect 2503 2144 2519 2208
rect 2583 2144 2599 2208
rect 2663 2144 2669 2208
rect 2353 2143 2669 2144
rect 3848 2208 4164 2209
rect 3848 2144 3854 2208
rect 3918 2144 3934 2208
rect 3998 2144 4014 2208
rect 4078 2144 4094 2208
rect 4158 2144 4164 2208
rect 3848 2143 4164 2144
rect 5343 2208 5659 2209
rect 5343 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5589 2208
rect 5653 2144 5659 2208
rect 5343 2143 5659 2144
rect 6838 2208 7154 2209
rect 6838 2144 6844 2208
rect 6908 2144 6924 2208
rect 6988 2144 7004 2208
rect 7068 2144 7084 2208
rect 7148 2144 7154 2208
rect 6838 2143 7154 2144
rect 7189 778 7255 781
rect 7411 778 8211 808
rect 7189 776 8211 778
rect 7189 720 7194 776
rect 7250 720 8211 776
rect 7189 718 8211 720
rect 7189 715 7255 718
rect 7411 688 8211 718
<< via3 >>
rect 1699 8188 1763 8192
rect 1699 8132 1703 8188
rect 1703 8132 1759 8188
rect 1759 8132 1763 8188
rect 1699 8128 1763 8132
rect 1779 8188 1843 8192
rect 1779 8132 1783 8188
rect 1783 8132 1839 8188
rect 1839 8132 1843 8188
rect 1779 8128 1843 8132
rect 1859 8188 1923 8192
rect 1859 8132 1863 8188
rect 1863 8132 1919 8188
rect 1919 8132 1923 8188
rect 1859 8128 1923 8132
rect 1939 8188 2003 8192
rect 1939 8132 1943 8188
rect 1943 8132 1999 8188
rect 1999 8132 2003 8188
rect 1939 8128 2003 8132
rect 3194 8188 3258 8192
rect 3194 8132 3198 8188
rect 3198 8132 3254 8188
rect 3254 8132 3258 8188
rect 3194 8128 3258 8132
rect 3274 8188 3338 8192
rect 3274 8132 3278 8188
rect 3278 8132 3334 8188
rect 3334 8132 3338 8188
rect 3274 8128 3338 8132
rect 3354 8188 3418 8192
rect 3354 8132 3358 8188
rect 3358 8132 3414 8188
rect 3414 8132 3418 8188
rect 3354 8128 3418 8132
rect 3434 8188 3498 8192
rect 3434 8132 3438 8188
rect 3438 8132 3494 8188
rect 3494 8132 3498 8188
rect 3434 8128 3498 8132
rect 4689 8188 4753 8192
rect 4689 8132 4693 8188
rect 4693 8132 4749 8188
rect 4749 8132 4753 8188
rect 4689 8128 4753 8132
rect 4769 8188 4833 8192
rect 4769 8132 4773 8188
rect 4773 8132 4829 8188
rect 4829 8132 4833 8188
rect 4769 8128 4833 8132
rect 4849 8188 4913 8192
rect 4849 8132 4853 8188
rect 4853 8132 4909 8188
rect 4909 8132 4913 8188
rect 4849 8128 4913 8132
rect 4929 8188 4993 8192
rect 4929 8132 4933 8188
rect 4933 8132 4989 8188
rect 4989 8132 4993 8188
rect 4929 8128 4993 8132
rect 6184 8188 6248 8192
rect 6184 8132 6188 8188
rect 6188 8132 6244 8188
rect 6244 8132 6248 8188
rect 6184 8128 6248 8132
rect 6264 8188 6328 8192
rect 6264 8132 6268 8188
rect 6268 8132 6324 8188
rect 6324 8132 6328 8188
rect 6264 8128 6328 8132
rect 6344 8188 6408 8192
rect 6344 8132 6348 8188
rect 6348 8132 6404 8188
rect 6404 8132 6408 8188
rect 6344 8128 6408 8132
rect 6424 8188 6488 8192
rect 6424 8132 6428 8188
rect 6428 8132 6484 8188
rect 6484 8132 6488 8188
rect 6424 8128 6488 8132
rect 2359 7644 2423 7648
rect 2359 7588 2363 7644
rect 2363 7588 2419 7644
rect 2419 7588 2423 7644
rect 2359 7584 2423 7588
rect 2439 7644 2503 7648
rect 2439 7588 2443 7644
rect 2443 7588 2499 7644
rect 2499 7588 2503 7644
rect 2439 7584 2503 7588
rect 2519 7644 2583 7648
rect 2519 7588 2523 7644
rect 2523 7588 2579 7644
rect 2579 7588 2583 7644
rect 2519 7584 2583 7588
rect 2599 7644 2663 7648
rect 2599 7588 2603 7644
rect 2603 7588 2659 7644
rect 2659 7588 2663 7644
rect 2599 7584 2663 7588
rect 3854 7644 3918 7648
rect 3854 7588 3858 7644
rect 3858 7588 3914 7644
rect 3914 7588 3918 7644
rect 3854 7584 3918 7588
rect 3934 7644 3998 7648
rect 3934 7588 3938 7644
rect 3938 7588 3994 7644
rect 3994 7588 3998 7644
rect 3934 7584 3998 7588
rect 4014 7644 4078 7648
rect 4014 7588 4018 7644
rect 4018 7588 4074 7644
rect 4074 7588 4078 7644
rect 4014 7584 4078 7588
rect 4094 7644 4158 7648
rect 4094 7588 4098 7644
rect 4098 7588 4154 7644
rect 4154 7588 4158 7644
rect 4094 7584 4158 7588
rect 5349 7644 5413 7648
rect 5349 7588 5353 7644
rect 5353 7588 5409 7644
rect 5409 7588 5413 7644
rect 5349 7584 5413 7588
rect 5429 7644 5493 7648
rect 5429 7588 5433 7644
rect 5433 7588 5489 7644
rect 5489 7588 5493 7644
rect 5429 7584 5493 7588
rect 5509 7644 5573 7648
rect 5509 7588 5513 7644
rect 5513 7588 5569 7644
rect 5569 7588 5573 7644
rect 5509 7584 5573 7588
rect 5589 7644 5653 7648
rect 5589 7588 5593 7644
rect 5593 7588 5649 7644
rect 5649 7588 5653 7644
rect 5589 7584 5653 7588
rect 6844 7644 6908 7648
rect 6844 7588 6848 7644
rect 6848 7588 6904 7644
rect 6904 7588 6908 7644
rect 6844 7584 6908 7588
rect 6924 7644 6988 7648
rect 6924 7588 6928 7644
rect 6928 7588 6984 7644
rect 6984 7588 6988 7644
rect 6924 7584 6988 7588
rect 7004 7644 7068 7648
rect 7004 7588 7008 7644
rect 7008 7588 7064 7644
rect 7064 7588 7068 7644
rect 7004 7584 7068 7588
rect 7084 7644 7148 7648
rect 7084 7588 7088 7644
rect 7088 7588 7144 7644
rect 7144 7588 7148 7644
rect 7084 7584 7148 7588
rect 1699 7100 1763 7104
rect 1699 7044 1703 7100
rect 1703 7044 1759 7100
rect 1759 7044 1763 7100
rect 1699 7040 1763 7044
rect 1779 7100 1843 7104
rect 1779 7044 1783 7100
rect 1783 7044 1839 7100
rect 1839 7044 1843 7100
rect 1779 7040 1843 7044
rect 1859 7100 1923 7104
rect 1859 7044 1863 7100
rect 1863 7044 1919 7100
rect 1919 7044 1923 7100
rect 1859 7040 1923 7044
rect 1939 7100 2003 7104
rect 1939 7044 1943 7100
rect 1943 7044 1999 7100
rect 1999 7044 2003 7100
rect 1939 7040 2003 7044
rect 3194 7100 3258 7104
rect 3194 7044 3198 7100
rect 3198 7044 3254 7100
rect 3254 7044 3258 7100
rect 3194 7040 3258 7044
rect 3274 7100 3338 7104
rect 3274 7044 3278 7100
rect 3278 7044 3334 7100
rect 3334 7044 3338 7100
rect 3274 7040 3338 7044
rect 3354 7100 3418 7104
rect 3354 7044 3358 7100
rect 3358 7044 3414 7100
rect 3414 7044 3418 7100
rect 3354 7040 3418 7044
rect 3434 7100 3498 7104
rect 3434 7044 3438 7100
rect 3438 7044 3494 7100
rect 3494 7044 3498 7100
rect 3434 7040 3498 7044
rect 4689 7100 4753 7104
rect 4689 7044 4693 7100
rect 4693 7044 4749 7100
rect 4749 7044 4753 7100
rect 4689 7040 4753 7044
rect 4769 7100 4833 7104
rect 4769 7044 4773 7100
rect 4773 7044 4829 7100
rect 4829 7044 4833 7100
rect 4769 7040 4833 7044
rect 4849 7100 4913 7104
rect 4849 7044 4853 7100
rect 4853 7044 4909 7100
rect 4909 7044 4913 7100
rect 4849 7040 4913 7044
rect 4929 7100 4993 7104
rect 4929 7044 4933 7100
rect 4933 7044 4989 7100
rect 4989 7044 4993 7100
rect 4929 7040 4993 7044
rect 6184 7100 6248 7104
rect 6184 7044 6188 7100
rect 6188 7044 6244 7100
rect 6244 7044 6248 7100
rect 6184 7040 6248 7044
rect 6264 7100 6328 7104
rect 6264 7044 6268 7100
rect 6268 7044 6324 7100
rect 6324 7044 6328 7100
rect 6264 7040 6328 7044
rect 6344 7100 6408 7104
rect 6344 7044 6348 7100
rect 6348 7044 6404 7100
rect 6404 7044 6408 7100
rect 6344 7040 6408 7044
rect 6424 7100 6488 7104
rect 6424 7044 6428 7100
rect 6428 7044 6484 7100
rect 6484 7044 6488 7100
rect 6424 7040 6488 7044
rect 2359 6556 2423 6560
rect 2359 6500 2363 6556
rect 2363 6500 2419 6556
rect 2419 6500 2423 6556
rect 2359 6496 2423 6500
rect 2439 6556 2503 6560
rect 2439 6500 2443 6556
rect 2443 6500 2499 6556
rect 2499 6500 2503 6556
rect 2439 6496 2503 6500
rect 2519 6556 2583 6560
rect 2519 6500 2523 6556
rect 2523 6500 2579 6556
rect 2579 6500 2583 6556
rect 2519 6496 2583 6500
rect 2599 6556 2663 6560
rect 2599 6500 2603 6556
rect 2603 6500 2659 6556
rect 2659 6500 2663 6556
rect 2599 6496 2663 6500
rect 3854 6556 3918 6560
rect 3854 6500 3858 6556
rect 3858 6500 3914 6556
rect 3914 6500 3918 6556
rect 3854 6496 3918 6500
rect 3934 6556 3998 6560
rect 3934 6500 3938 6556
rect 3938 6500 3994 6556
rect 3994 6500 3998 6556
rect 3934 6496 3998 6500
rect 4014 6556 4078 6560
rect 4014 6500 4018 6556
rect 4018 6500 4074 6556
rect 4074 6500 4078 6556
rect 4014 6496 4078 6500
rect 4094 6556 4158 6560
rect 4094 6500 4098 6556
rect 4098 6500 4154 6556
rect 4154 6500 4158 6556
rect 4094 6496 4158 6500
rect 5349 6556 5413 6560
rect 5349 6500 5353 6556
rect 5353 6500 5409 6556
rect 5409 6500 5413 6556
rect 5349 6496 5413 6500
rect 5429 6556 5493 6560
rect 5429 6500 5433 6556
rect 5433 6500 5489 6556
rect 5489 6500 5493 6556
rect 5429 6496 5493 6500
rect 5509 6556 5573 6560
rect 5509 6500 5513 6556
rect 5513 6500 5569 6556
rect 5569 6500 5573 6556
rect 5509 6496 5573 6500
rect 5589 6556 5653 6560
rect 5589 6500 5593 6556
rect 5593 6500 5649 6556
rect 5649 6500 5653 6556
rect 5589 6496 5653 6500
rect 6844 6556 6908 6560
rect 6844 6500 6848 6556
rect 6848 6500 6904 6556
rect 6904 6500 6908 6556
rect 6844 6496 6908 6500
rect 6924 6556 6988 6560
rect 6924 6500 6928 6556
rect 6928 6500 6984 6556
rect 6984 6500 6988 6556
rect 6924 6496 6988 6500
rect 7004 6556 7068 6560
rect 7004 6500 7008 6556
rect 7008 6500 7064 6556
rect 7064 6500 7068 6556
rect 7004 6496 7068 6500
rect 7084 6556 7148 6560
rect 7084 6500 7088 6556
rect 7088 6500 7144 6556
rect 7144 6500 7148 6556
rect 7084 6496 7148 6500
rect 1699 6012 1763 6016
rect 1699 5956 1703 6012
rect 1703 5956 1759 6012
rect 1759 5956 1763 6012
rect 1699 5952 1763 5956
rect 1779 6012 1843 6016
rect 1779 5956 1783 6012
rect 1783 5956 1839 6012
rect 1839 5956 1843 6012
rect 1779 5952 1843 5956
rect 1859 6012 1923 6016
rect 1859 5956 1863 6012
rect 1863 5956 1919 6012
rect 1919 5956 1923 6012
rect 1859 5952 1923 5956
rect 1939 6012 2003 6016
rect 1939 5956 1943 6012
rect 1943 5956 1999 6012
rect 1999 5956 2003 6012
rect 1939 5952 2003 5956
rect 3194 6012 3258 6016
rect 3194 5956 3198 6012
rect 3198 5956 3254 6012
rect 3254 5956 3258 6012
rect 3194 5952 3258 5956
rect 3274 6012 3338 6016
rect 3274 5956 3278 6012
rect 3278 5956 3334 6012
rect 3334 5956 3338 6012
rect 3274 5952 3338 5956
rect 3354 6012 3418 6016
rect 3354 5956 3358 6012
rect 3358 5956 3414 6012
rect 3414 5956 3418 6012
rect 3354 5952 3418 5956
rect 3434 6012 3498 6016
rect 3434 5956 3438 6012
rect 3438 5956 3494 6012
rect 3494 5956 3498 6012
rect 3434 5952 3498 5956
rect 4689 6012 4753 6016
rect 4689 5956 4693 6012
rect 4693 5956 4749 6012
rect 4749 5956 4753 6012
rect 4689 5952 4753 5956
rect 4769 6012 4833 6016
rect 4769 5956 4773 6012
rect 4773 5956 4829 6012
rect 4829 5956 4833 6012
rect 4769 5952 4833 5956
rect 4849 6012 4913 6016
rect 4849 5956 4853 6012
rect 4853 5956 4909 6012
rect 4909 5956 4913 6012
rect 4849 5952 4913 5956
rect 4929 6012 4993 6016
rect 4929 5956 4933 6012
rect 4933 5956 4989 6012
rect 4989 5956 4993 6012
rect 4929 5952 4993 5956
rect 6184 6012 6248 6016
rect 6184 5956 6188 6012
rect 6188 5956 6244 6012
rect 6244 5956 6248 6012
rect 6184 5952 6248 5956
rect 6264 6012 6328 6016
rect 6264 5956 6268 6012
rect 6268 5956 6324 6012
rect 6324 5956 6328 6012
rect 6264 5952 6328 5956
rect 6344 6012 6408 6016
rect 6344 5956 6348 6012
rect 6348 5956 6404 6012
rect 6404 5956 6408 6012
rect 6344 5952 6408 5956
rect 6424 6012 6488 6016
rect 6424 5956 6428 6012
rect 6428 5956 6484 6012
rect 6484 5956 6488 6012
rect 6424 5952 6488 5956
rect 2359 5468 2423 5472
rect 2359 5412 2363 5468
rect 2363 5412 2419 5468
rect 2419 5412 2423 5468
rect 2359 5408 2423 5412
rect 2439 5468 2503 5472
rect 2439 5412 2443 5468
rect 2443 5412 2499 5468
rect 2499 5412 2503 5468
rect 2439 5408 2503 5412
rect 2519 5468 2583 5472
rect 2519 5412 2523 5468
rect 2523 5412 2579 5468
rect 2579 5412 2583 5468
rect 2519 5408 2583 5412
rect 2599 5468 2663 5472
rect 2599 5412 2603 5468
rect 2603 5412 2659 5468
rect 2659 5412 2663 5468
rect 2599 5408 2663 5412
rect 3854 5468 3918 5472
rect 3854 5412 3858 5468
rect 3858 5412 3914 5468
rect 3914 5412 3918 5468
rect 3854 5408 3918 5412
rect 3934 5468 3998 5472
rect 3934 5412 3938 5468
rect 3938 5412 3994 5468
rect 3994 5412 3998 5468
rect 3934 5408 3998 5412
rect 4014 5468 4078 5472
rect 4014 5412 4018 5468
rect 4018 5412 4074 5468
rect 4074 5412 4078 5468
rect 4014 5408 4078 5412
rect 4094 5468 4158 5472
rect 4094 5412 4098 5468
rect 4098 5412 4154 5468
rect 4154 5412 4158 5468
rect 4094 5408 4158 5412
rect 5349 5468 5413 5472
rect 5349 5412 5353 5468
rect 5353 5412 5409 5468
rect 5409 5412 5413 5468
rect 5349 5408 5413 5412
rect 5429 5468 5493 5472
rect 5429 5412 5433 5468
rect 5433 5412 5489 5468
rect 5489 5412 5493 5468
rect 5429 5408 5493 5412
rect 5509 5468 5573 5472
rect 5509 5412 5513 5468
rect 5513 5412 5569 5468
rect 5569 5412 5573 5468
rect 5509 5408 5573 5412
rect 5589 5468 5653 5472
rect 5589 5412 5593 5468
rect 5593 5412 5649 5468
rect 5649 5412 5653 5468
rect 5589 5408 5653 5412
rect 6844 5468 6908 5472
rect 6844 5412 6848 5468
rect 6848 5412 6904 5468
rect 6904 5412 6908 5468
rect 6844 5408 6908 5412
rect 6924 5468 6988 5472
rect 6924 5412 6928 5468
rect 6928 5412 6984 5468
rect 6984 5412 6988 5468
rect 6924 5408 6988 5412
rect 7004 5468 7068 5472
rect 7004 5412 7008 5468
rect 7008 5412 7064 5468
rect 7064 5412 7068 5468
rect 7004 5408 7068 5412
rect 7084 5468 7148 5472
rect 7084 5412 7088 5468
rect 7088 5412 7144 5468
rect 7144 5412 7148 5468
rect 7084 5408 7148 5412
rect 1699 4924 1763 4928
rect 1699 4868 1703 4924
rect 1703 4868 1759 4924
rect 1759 4868 1763 4924
rect 1699 4864 1763 4868
rect 1779 4924 1843 4928
rect 1779 4868 1783 4924
rect 1783 4868 1839 4924
rect 1839 4868 1843 4924
rect 1779 4864 1843 4868
rect 1859 4924 1923 4928
rect 1859 4868 1863 4924
rect 1863 4868 1919 4924
rect 1919 4868 1923 4924
rect 1859 4864 1923 4868
rect 1939 4924 2003 4928
rect 1939 4868 1943 4924
rect 1943 4868 1999 4924
rect 1999 4868 2003 4924
rect 1939 4864 2003 4868
rect 3194 4924 3258 4928
rect 3194 4868 3198 4924
rect 3198 4868 3254 4924
rect 3254 4868 3258 4924
rect 3194 4864 3258 4868
rect 3274 4924 3338 4928
rect 3274 4868 3278 4924
rect 3278 4868 3334 4924
rect 3334 4868 3338 4924
rect 3274 4864 3338 4868
rect 3354 4924 3418 4928
rect 3354 4868 3358 4924
rect 3358 4868 3414 4924
rect 3414 4868 3418 4924
rect 3354 4864 3418 4868
rect 3434 4924 3498 4928
rect 3434 4868 3438 4924
rect 3438 4868 3494 4924
rect 3494 4868 3498 4924
rect 3434 4864 3498 4868
rect 4689 4924 4753 4928
rect 4689 4868 4693 4924
rect 4693 4868 4749 4924
rect 4749 4868 4753 4924
rect 4689 4864 4753 4868
rect 4769 4924 4833 4928
rect 4769 4868 4773 4924
rect 4773 4868 4829 4924
rect 4829 4868 4833 4924
rect 4769 4864 4833 4868
rect 4849 4924 4913 4928
rect 4849 4868 4853 4924
rect 4853 4868 4909 4924
rect 4909 4868 4913 4924
rect 4849 4864 4913 4868
rect 4929 4924 4993 4928
rect 4929 4868 4933 4924
rect 4933 4868 4989 4924
rect 4989 4868 4993 4924
rect 4929 4864 4993 4868
rect 6184 4924 6248 4928
rect 6184 4868 6188 4924
rect 6188 4868 6244 4924
rect 6244 4868 6248 4924
rect 6184 4864 6248 4868
rect 6264 4924 6328 4928
rect 6264 4868 6268 4924
rect 6268 4868 6324 4924
rect 6324 4868 6328 4924
rect 6264 4864 6328 4868
rect 6344 4924 6408 4928
rect 6344 4868 6348 4924
rect 6348 4868 6404 4924
rect 6404 4868 6408 4924
rect 6344 4864 6408 4868
rect 6424 4924 6488 4928
rect 6424 4868 6428 4924
rect 6428 4868 6484 4924
rect 6484 4868 6488 4924
rect 6424 4864 6488 4868
rect 2359 4380 2423 4384
rect 2359 4324 2363 4380
rect 2363 4324 2419 4380
rect 2419 4324 2423 4380
rect 2359 4320 2423 4324
rect 2439 4380 2503 4384
rect 2439 4324 2443 4380
rect 2443 4324 2499 4380
rect 2499 4324 2503 4380
rect 2439 4320 2503 4324
rect 2519 4380 2583 4384
rect 2519 4324 2523 4380
rect 2523 4324 2579 4380
rect 2579 4324 2583 4380
rect 2519 4320 2583 4324
rect 2599 4380 2663 4384
rect 2599 4324 2603 4380
rect 2603 4324 2659 4380
rect 2659 4324 2663 4380
rect 2599 4320 2663 4324
rect 3854 4380 3918 4384
rect 3854 4324 3858 4380
rect 3858 4324 3914 4380
rect 3914 4324 3918 4380
rect 3854 4320 3918 4324
rect 3934 4380 3998 4384
rect 3934 4324 3938 4380
rect 3938 4324 3994 4380
rect 3994 4324 3998 4380
rect 3934 4320 3998 4324
rect 4014 4380 4078 4384
rect 4014 4324 4018 4380
rect 4018 4324 4074 4380
rect 4074 4324 4078 4380
rect 4014 4320 4078 4324
rect 4094 4380 4158 4384
rect 4094 4324 4098 4380
rect 4098 4324 4154 4380
rect 4154 4324 4158 4380
rect 4094 4320 4158 4324
rect 5349 4380 5413 4384
rect 5349 4324 5353 4380
rect 5353 4324 5409 4380
rect 5409 4324 5413 4380
rect 5349 4320 5413 4324
rect 5429 4380 5493 4384
rect 5429 4324 5433 4380
rect 5433 4324 5489 4380
rect 5489 4324 5493 4380
rect 5429 4320 5493 4324
rect 5509 4380 5573 4384
rect 5509 4324 5513 4380
rect 5513 4324 5569 4380
rect 5569 4324 5573 4380
rect 5509 4320 5573 4324
rect 5589 4380 5653 4384
rect 5589 4324 5593 4380
rect 5593 4324 5649 4380
rect 5649 4324 5653 4380
rect 5589 4320 5653 4324
rect 6844 4380 6908 4384
rect 6844 4324 6848 4380
rect 6848 4324 6904 4380
rect 6904 4324 6908 4380
rect 6844 4320 6908 4324
rect 6924 4380 6988 4384
rect 6924 4324 6928 4380
rect 6928 4324 6984 4380
rect 6984 4324 6988 4380
rect 6924 4320 6988 4324
rect 7004 4380 7068 4384
rect 7004 4324 7008 4380
rect 7008 4324 7064 4380
rect 7064 4324 7068 4380
rect 7004 4320 7068 4324
rect 7084 4380 7148 4384
rect 7084 4324 7088 4380
rect 7088 4324 7144 4380
rect 7144 4324 7148 4380
rect 7084 4320 7148 4324
rect 1699 3836 1763 3840
rect 1699 3780 1703 3836
rect 1703 3780 1759 3836
rect 1759 3780 1763 3836
rect 1699 3776 1763 3780
rect 1779 3836 1843 3840
rect 1779 3780 1783 3836
rect 1783 3780 1839 3836
rect 1839 3780 1843 3836
rect 1779 3776 1843 3780
rect 1859 3836 1923 3840
rect 1859 3780 1863 3836
rect 1863 3780 1919 3836
rect 1919 3780 1923 3836
rect 1859 3776 1923 3780
rect 1939 3836 2003 3840
rect 1939 3780 1943 3836
rect 1943 3780 1999 3836
rect 1999 3780 2003 3836
rect 1939 3776 2003 3780
rect 3194 3836 3258 3840
rect 3194 3780 3198 3836
rect 3198 3780 3254 3836
rect 3254 3780 3258 3836
rect 3194 3776 3258 3780
rect 3274 3836 3338 3840
rect 3274 3780 3278 3836
rect 3278 3780 3334 3836
rect 3334 3780 3338 3836
rect 3274 3776 3338 3780
rect 3354 3836 3418 3840
rect 3354 3780 3358 3836
rect 3358 3780 3414 3836
rect 3414 3780 3418 3836
rect 3354 3776 3418 3780
rect 3434 3836 3498 3840
rect 3434 3780 3438 3836
rect 3438 3780 3494 3836
rect 3494 3780 3498 3836
rect 3434 3776 3498 3780
rect 4689 3836 4753 3840
rect 4689 3780 4693 3836
rect 4693 3780 4749 3836
rect 4749 3780 4753 3836
rect 4689 3776 4753 3780
rect 4769 3836 4833 3840
rect 4769 3780 4773 3836
rect 4773 3780 4829 3836
rect 4829 3780 4833 3836
rect 4769 3776 4833 3780
rect 4849 3836 4913 3840
rect 4849 3780 4853 3836
rect 4853 3780 4909 3836
rect 4909 3780 4913 3836
rect 4849 3776 4913 3780
rect 4929 3836 4993 3840
rect 4929 3780 4933 3836
rect 4933 3780 4989 3836
rect 4989 3780 4993 3836
rect 4929 3776 4993 3780
rect 6184 3836 6248 3840
rect 6184 3780 6188 3836
rect 6188 3780 6244 3836
rect 6244 3780 6248 3836
rect 6184 3776 6248 3780
rect 6264 3836 6328 3840
rect 6264 3780 6268 3836
rect 6268 3780 6324 3836
rect 6324 3780 6328 3836
rect 6264 3776 6328 3780
rect 6344 3836 6408 3840
rect 6344 3780 6348 3836
rect 6348 3780 6404 3836
rect 6404 3780 6408 3836
rect 6344 3776 6408 3780
rect 6424 3836 6488 3840
rect 6424 3780 6428 3836
rect 6428 3780 6484 3836
rect 6484 3780 6488 3836
rect 6424 3776 6488 3780
rect 2359 3292 2423 3296
rect 2359 3236 2363 3292
rect 2363 3236 2419 3292
rect 2419 3236 2423 3292
rect 2359 3232 2423 3236
rect 2439 3292 2503 3296
rect 2439 3236 2443 3292
rect 2443 3236 2499 3292
rect 2499 3236 2503 3292
rect 2439 3232 2503 3236
rect 2519 3292 2583 3296
rect 2519 3236 2523 3292
rect 2523 3236 2579 3292
rect 2579 3236 2583 3292
rect 2519 3232 2583 3236
rect 2599 3292 2663 3296
rect 2599 3236 2603 3292
rect 2603 3236 2659 3292
rect 2659 3236 2663 3292
rect 2599 3232 2663 3236
rect 3854 3292 3918 3296
rect 3854 3236 3858 3292
rect 3858 3236 3914 3292
rect 3914 3236 3918 3292
rect 3854 3232 3918 3236
rect 3934 3292 3998 3296
rect 3934 3236 3938 3292
rect 3938 3236 3994 3292
rect 3994 3236 3998 3292
rect 3934 3232 3998 3236
rect 4014 3292 4078 3296
rect 4014 3236 4018 3292
rect 4018 3236 4074 3292
rect 4074 3236 4078 3292
rect 4014 3232 4078 3236
rect 4094 3292 4158 3296
rect 4094 3236 4098 3292
rect 4098 3236 4154 3292
rect 4154 3236 4158 3292
rect 4094 3232 4158 3236
rect 5349 3292 5413 3296
rect 5349 3236 5353 3292
rect 5353 3236 5409 3292
rect 5409 3236 5413 3292
rect 5349 3232 5413 3236
rect 5429 3292 5493 3296
rect 5429 3236 5433 3292
rect 5433 3236 5489 3292
rect 5489 3236 5493 3292
rect 5429 3232 5493 3236
rect 5509 3292 5573 3296
rect 5509 3236 5513 3292
rect 5513 3236 5569 3292
rect 5569 3236 5573 3292
rect 5509 3232 5573 3236
rect 5589 3292 5653 3296
rect 5589 3236 5593 3292
rect 5593 3236 5649 3292
rect 5649 3236 5653 3292
rect 5589 3232 5653 3236
rect 6844 3292 6908 3296
rect 6844 3236 6848 3292
rect 6848 3236 6904 3292
rect 6904 3236 6908 3292
rect 6844 3232 6908 3236
rect 6924 3292 6988 3296
rect 6924 3236 6928 3292
rect 6928 3236 6984 3292
rect 6984 3236 6988 3292
rect 6924 3232 6988 3236
rect 7004 3292 7068 3296
rect 7004 3236 7008 3292
rect 7008 3236 7064 3292
rect 7064 3236 7068 3292
rect 7004 3232 7068 3236
rect 7084 3292 7148 3296
rect 7084 3236 7088 3292
rect 7088 3236 7144 3292
rect 7144 3236 7148 3292
rect 7084 3232 7148 3236
rect 1699 2748 1763 2752
rect 1699 2692 1703 2748
rect 1703 2692 1759 2748
rect 1759 2692 1763 2748
rect 1699 2688 1763 2692
rect 1779 2748 1843 2752
rect 1779 2692 1783 2748
rect 1783 2692 1839 2748
rect 1839 2692 1843 2748
rect 1779 2688 1843 2692
rect 1859 2748 1923 2752
rect 1859 2692 1863 2748
rect 1863 2692 1919 2748
rect 1919 2692 1923 2748
rect 1859 2688 1923 2692
rect 1939 2748 2003 2752
rect 1939 2692 1943 2748
rect 1943 2692 1999 2748
rect 1999 2692 2003 2748
rect 1939 2688 2003 2692
rect 3194 2748 3258 2752
rect 3194 2692 3198 2748
rect 3198 2692 3254 2748
rect 3254 2692 3258 2748
rect 3194 2688 3258 2692
rect 3274 2748 3338 2752
rect 3274 2692 3278 2748
rect 3278 2692 3334 2748
rect 3334 2692 3338 2748
rect 3274 2688 3338 2692
rect 3354 2748 3418 2752
rect 3354 2692 3358 2748
rect 3358 2692 3414 2748
rect 3414 2692 3418 2748
rect 3354 2688 3418 2692
rect 3434 2748 3498 2752
rect 3434 2692 3438 2748
rect 3438 2692 3494 2748
rect 3494 2692 3498 2748
rect 3434 2688 3498 2692
rect 4689 2748 4753 2752
rect 4689 2692 4693 2748
rect 4693 2692 4749 2748
rect 4749 2692 4753 2748
rect 4689 2688 4753 2692
rect 4769 2748 4833 2752
rect 4769 2692 4773 2748
rect 4773 2692 4829 2748
rect 4829 2692 4833 2748
rect 4769 2688 4833 2692
rect 4849 2748 4913 2752
rect 4849 2692 4853 2748
rect 4853 2692 4909 2748
rect 4909 2692 4913 2748
rect 4849 2688 4913 2692
rect 4929 2748 4993 2752
rect 4929 2692 4933 2748
rect 4933 2692 4989 2748
rect 4989 2692 4993 2748
rect 4929 2688 4993 2692
rect 6184 2748 6248 2752
rect 6184 2692 6188 2748
rect 6188 2692 6244 2748
rect 6244 2692 6248 2748
rect 6184 2688 6248 2692
rect 6264 2748 6328 2752
rect 6264 2692 6268 2748
rect 6268 2692 6324 2748
rect 6324 2692 6328 2748
rect 6264 2688 6328 2692
rect 6344 2748 6408 2752
rect 6344 2692 6348 2748
rect 6348 2692 6404 2748
rect 6404 2692 6408 2748
rect 6344 2688 6408 2692
rect 6424 2748 6488 2752
rect 6424 2692 6428 2748
rect 6428 2692 6484 2748
rect 6484 2692 6488 2748
rect 6424 2688 6488 2692
rect 2359 2204 2423 2208
rect 2359 2148 2363 2204
rect 2363 2148 2419 2204
rect 2419 2148 2423 2204
rect 2359 2144 2423 2148
rect 2439 2204 2503 2208
rect 2439 2148 2443 2204
rect 2443 2148 2499 2204
rect 2499 2148 2503 2204
rect 2439 2144 2503 2148
rect 2519 2204 2583 2208
rect 2519 2148 2523 2204
rect 2523 2148 2579 2204
rect 2579 2148 2583 2204
rect 2519 2144 2583 2148
rect 2599 2204 2663 2208
rect 2599 2148 2603 2204
rect 2603 2148 2659 2204
rect 2659 2148 2663 2204
rect 2599 2144 2663 2148
rect 3854 2204 3918 2208
rect 3854 2148 3858 2204
rect 3858 2148 3914 2204
rect 3914 2148 3918 2204
rect 3854 2144 3918 2148
rect 3934 2204 3998 2208
rect 3934 2148 3938 2204
rect 3938 2148 3994 2204
rect 3994 2148 3998 2204
rect 3934 2144 3998 2148
rect 4014 2204 4078 2208
rect 4014 2148 4018 2204
rect 4018 2148 4074 2204
rect 4074 2148 4078 2204
rect 4014 2144 4078 2148
rect 4094 2204 4158 2208
rect 4094 2148 4098 2204
rect 4098 2148 4154 2204
rect 4154 2148 4158 2204
rect 4094 2144 4158 2148
rect 5349 2204 5413 2208
rect 5349 2148 5353 2204
rect 5353 2148 5409 2204
rect 5409 2148 5413 2204
rect 5349 2144 5413 2148
rect 5429 2204 5493 2208
rect 5429 2148 5433 2204
rect 5433 2148 5489 2204
rect 5489 2148 5493 2204
rect 5429 2144 5493 2148
rect 5509 2204 5573 2208
rect 5509 2148 5513 2204
rect 5513 2148 5569 2204
rect 5569 2148 5573 2204
rect 5509 2144 5573 2148
rect 5589 2204 5653 2208
rect 5589 2148 5593 2204
rect 5593 2148 5649 2204
rect 5649 2148 5653 2204
rect 5589 2144 5653 2148
rect 6844 2204 6908 2208
rect 6844 2148 6848 2204
rect 6848 2148 6904 2204
rect 6904 2148 6908 2204
rect 6844 2144 6908 2148
rect 6924 2204 6988 2208
rect 6924 2148 6928 2204
rect 6928 2148 6984 2204
rect 6984 2148 6988 2204
rect 6924 2144 6988 2148
rect 7004 2204 7068 2208
rect 7004 2148 7008 2204
rect 7008 2148 7064 2204
rect 7064 2148 7068 2204
rect 7004 2144 7068 2148
rect 7084 2204 7148 2208
rect 7084 2148 7088 2204
rect 7088 2148 7144 2204
rect 7144 2148 7148 2204
rect 7084 2144 7148 2148
<< metal4 >>
rect 1691 8192 2011 8208
rect 1691 8128 1699 8192
rect 1763 8128 1779 8192
rect 1843 8128 1859 8192
rect 1923 8128 1939 8192
rect 2003 8128 2011 8192
rect 1691 7526 2011 8128
rect 1691 7290 1733 7526
rect 1969 7290 2011 7526
rect 1691 7104 2011 7290
rect 1691 7040 1699 7104
rect 1763 7040 1779 7104
rect 1843 7040 1859 7104
rect 1923 7040 1939 7104
rect 2003 7040 2011 7104
rect 1691 6031 2011 7040
rect 1691 6016 1733 6031
rect 1969 6016 2011 6031
rect 1691 5952 1699 6016
rect 2003 5952 2011 6016
rect 1691 5795 1733 5952
rect 1969 5795 2011 5952
rect 1691 4928 2011 5795
rect 1691 4864 1699 4928
rect 1763 4864 1779 4928
rect 1843 4864 1859 4928
rect 1923 4864 1939 4928
rect 2003 4864 2011 4928
rect 1691 4536 2011 4864
rect 1691 4300 1733 4536
rect 1969 4300 2011 4536
rect 1691 3840 2011 4300
rect 1691 3776 1699 3840
rect 1763 3776 1779 3840
rect 1843 3776 1859 3840
rect 1923 3776 1939 3840
rect 2003 3776 2011 3840
rect 1691 3041 2011 3776
rect 1691 2805 1733 3041
rect 1969 2805 2011 3041
rect 1691 2752 2011 2805
rect 1691 2688 1699 2752
rect 1763 2688 1779 2752
rect 1843 2688 1859 2752
rect 1923 2688 1939 2752
rect 2003 2688 2011 2752
rect 1691 2128 2011 2688
rect 2351 8186 2671 8228
rect 2351 7950 2393 8186
rect 2629 7950 2671 8186
rect 2351 7648 2671 7950
rect 2351 7584 2359 7648
rect 2423 7584 2439 7648
rect 2503 7584 2519 7648
rect 2583 7584 2599 7648
rect 2663 7584 2671 7648
rect 2351 6691 2671 7584
rect 2351 6560 2393 6691
rect 2629 6560 2671 6691
rect 2351 6496 2359 6560
rect 2663 6496 2671 6560
rect 2351 6455 2393 6496
rect 2629 6455 2671 6496
rect 2351 5472 2671 6455
rect 2351 5408 2359 5472
rect 2423 5408 2439 5472
rect 2503 5408 2519 5472
rect 2583 5408 2599 5472
rect 2663 5408 2671 5472
rect 2351 5196 2671 5408
rect 2351 4960 2393 5196
rect 2629 4960 2671 5196
rect 2351 4384 2671 4960
rect 2351 4320 2359 4384
rect 2423 4320 2439 4384
rect 2503 4320 2519 4384
rect 2583 4320 2599 4384
rect 2663 4320 2671 4384
rect 2351 3701 2671 4320
rect 2351 3465 2393 3701
rect 2629 3465 2671 3701
rect 2351 3296 2671 3465
rect 2351 3232 2359 3296
rect 2423 3232 2439 3296
rect 2503 3232 2519 3296
rect 2583 3232 2599 3296
rect 2663 3232 2671 3296
rect 2351 2208 2671 3232
rect 2351 2144 2359 2208
rect 2423 2144 2439 2208
rect 2503 2144 2519 2208
rect 2583 2144 2599 2208
rect 2663 2144 2671 2208
rect 2351 2128 2671 2144
rect 3186 8192 3506 8208
rect 3186 8128 3194 8192
rect 3258 8128 3274 8192
rect 3338 8128 3354 8192
rect 3418 8128 3434 8192
rect 3498 8128 3506 8192
rect 3186 7526 3506 8128
rect 3186 7290 3228 7526
rect 3464 7290 3506 7526
rect 3186 7104 3506 7290
rect 3186 7040 3194 7104
rect 3258 7040 3274 7104
rect 3338 7040 3354 7104
rect 3418 7040 3434 7104
rect 3498 7040 3506 7104
rect 3186 6031 3506 7040
rect 3186 6016 3228 6031
rect 3464 6016 3506 6031
rect 3186 5952 3194 6016
rect 3498 5952 3506 6016
rect 3186 5795 3228 5952
rect 3464 5795 3506 5952
rect 3186 4928 3506 5795
rect 3186 4864 3194 4928
rect 3258 4864 3274 4928
rect 3338 4864 3354 4928
rect 3418 4864 3434 4928
rect 3498 4864 3506 4928
rect 3186 4536 3506 4864
rect 3186 4300 3228 4536
rect 3464 4300 3506 4536
rect 3186 3840 3506 4300
rect 3186 3776 3194 3840
rect 3258 3776 3274 3840
rect 3338 3776 3354 3840
rect 3418 3776 3434 3840
rect 3498 3776 3506 3840
rect 3186 3041 3506 3776
rect 3186 2805 3228 3041
rect 3464 2805 3506 3041
rect 3186 2752 3506 2805
rect 3186 2688 3194 2752
rect 3258 2688 3274 2752
rect 3338 2688 3354 2752
rect 3418 2688 3434 2752
rect 3498 2688 3506 2752
rect 3186 2128 3506 2688
rect 3846 8186 4166 8228
rect 3846 7950 3888 8186
rect 4124 7950 4166 8186
rect 3846 7648 4166 7950
rect 3846 7584 3854 7648
rect 3918 7584 3934 7648
rect 3998 7584 4014 7648
rect 4078 7584 4094 7648
rect 4158 7584 4166 7648
rect 3846 6691 4166 7584
rect 3846 6560 3888 6691
rect 4124 6560 4166 6691
rect 3846 6496 3854 6560
rect 4158 6496 4166 6560
rect 3846 6455 3888 6496
rect 4124 6455 4166 6496
rect 3846 5472 4166 6455
rect 3846 5408 3854 5472
rect 3918 5408 3934 5472
rect 3998 5408 4014 5472
rect 4078 5408 4094 5472
rect 4158 5408 4166 5472
rect 3846 5196 4166 5408
rect 3846 4960 3888 5196
rect 4124 4960 4166 5196
rect 3846 4384 4166 4960
rect 3846 4320 3854 4384
rect 3918 4320 3934 4384
rect 3998 4320 4014 4384
rect 4078 4320 4094 4384
rect 4158 4320 4166 4384
rect 3846 3701 4166 4320
rect 3846 3465 3888 3701
rect 4124 3465 4166 3701
rect 3846 3296 4166 3465
rect 3846 3232 3854 3296
rect 3918 3232 3934 3296
rect 3998 3232 4014 3296
rect 4078 3232 4094 3296
rect 4158 3232 4166 3296
rect 3846 2208 4166 3232
rect 3846 2144 3854 2208
rect 3918 2144 3934 2208
rect 3998 2144 4014 2208
rect 4078 2144 4094 2208
rect 4158 2144 4166 2208
rect 3846 2128 4166 2144
rect 4681 8192 5001 8208
rect 4681 8128 4689 8192
rect 4753 8128 4769 8192
rect 4833 8128 4849 8192
rect 4913 8128 4929 8192
rect 4993 8128 5001 8192
rect 4681 7526 5001 8128
rect 4681 7290 4723 7526
rect 4959 7290 5001 7526
rect 4681 7104 5001 7290
rect 4681 7040 4689 7104
rect 4753 7040 4769 7104
rect 4833 7040 4849 7104
rect 4913 7040 4929 7104
rect 4993 7040 5001 7104
rect 4681 6031 5001 7040
rect 4681 6016 4723 6031
rect 4959 6016 5001 6031
rect 4681 5952 4689 6016
rect 4993 5952 5001 6016
rect 4681 5795 4723 5952
rect 4959 5795 5001 5952
rect 4681 4928 5001 5795
rect 4681 4864 4689 4928
rect 4753 4864 4769 4928
rect 4833 4864 4849 4928
rect 4913 4864 4929 4928
rect 4993 4864 5001 4928
rect 4681 4536 5001 4864
rect 4681 4300 4723 4536
rect 4959 4300 5001 4536
rect 4681 3840 5001 4300
rect 4681 3776 4689 3840
rect 4753 3776 4769 3840
rect 4833 3776 4849 3840
rect 4913 3776 4929 3840
rect 4993 3776 5001 3840
rect 4681 3041 5001 3776
rect 4681 2805 4723 3041
rect 4959 2805 5001 3041
rect 4681 2752 5001 2805
rect 4681 2688 4689 2752
rect 4753 2688 4769 2752
rect 4833 2688 4849 2752
rect 4913 2688 4929 2752
rect 4993 2688 5001 2752
rect 4681 2128 5001 2688
rect 5341 8186 5661 8228
rect 5341 7950 5383 8186
rect 5619 7950 5661 8186
rect 5341 7648 5661 7950
rect 5341 7584 5349 7648
rect 5413 7584 5429 7648
rect 5493 7584 5509 7648
rect 5573 7584 5589 7648
rect 5653 7584 5661 7648
rect 5341 6691 5661 7584
rect 5341 6560 5383 6691
rect 5619 6560 5661 6691
rect 5341 6496 5349 6560
rect 5653 6496 5661 6560
rect 5341 6455 5383 6496
rect 5619 6455 5661 6496
rect 5341 5472 5661 6455
rect 5341 5408 5349 5472
rect 5413 5408 5429 5472
rect 5493 5408 5509 5472
rect 5573 5408 5589 5472
rect 5653 5408 5661 5472
rect 5341 5196 5661 5408
rect 5341 4960 5383 5196
rect 5619 4960 5661 5196
rect 5341 4384 5661 4960
rect 5341 4320 5349 4384
rect 5413 4320 5429 4384
rect 5493 4320 5509 4384
rect 5573 4320 5589 4384
rect 5653 4320 5661 4384
rect 5341 3701 5661 4320
rect 5341 3465 5383 3701
rect 5619 3465 5661 3701
rect 5341 3296 5661 3465
rect 5341 3232 5349 3296
rect 5413 3232 5429 3296
rect 5493 3232 5509 3296
rect 5573 3232 5589 3296
rect 5653 3232 5661 3296
rect 5341 2208 5661 3232
rect 5341 2144 5349 2208
rect 5413 2144 5429 2208
rect 5493 2144 5509 2208
rect 5573 2144 5589 2208
rect 5653 2144 5661 2208
rect 5341 2128 5661 2144
rect 6176 8192 6496 8208
rect 6176 8128 6184 8192
rect 6248 8128 6264 8192
rect 6328 8128 6344 8192
rect 6408 8128 6424 8192
rect 6488 8128 6496 8192
rect 6176 7526 6496 8128
rect 6176 7290 6218 7526
rect 6454 7290 6496 7526
rect 6176 7104 6496 7290
rect 6176 7040 6184 7104
rect 6248 7040 6264 7104
rect 6328 7040 6344 7104
rect 6408 7040 6424 7104
rect 6488 7040 6496 7104
rect 6176 6031 6496 7040
rect 6176 6016 6218 6031
rect 6454 6016 6496 6031
rect 6176 5952 6184 6016
rect 6488 5952 6496 6016
rect 6176 5795 6218 5952
rect 6454 5795 6496 5952
rect 6176 4928 6496 5795
rect 6176 4864 6184 4928
rect 6248 4864 6264 4928
rect 6328 4864 6344 4928
rect 6408 4864 6424 4928
rect 6488 4864 6496 4928
rect 6176 4536 6496 4864
rect 6176 4300 6218 4536
rect 6454 4300 6496 4536
rect 6176 3840 6496 4300
rect 6176 3776 6184 3840
rect 6248 3776 6264 3840
rect 6328 3776 6344 3840
rect 6408 3776 6424 3840
rect 6488 3776 6496 3840
rect 6176 3041 6496 3776
rect 6176 2805 6218 3041
rect 6454 2805 6496 3041
rect 6176 2752 6496 2805
rect 6176 2688 6184 2752
rect 6248 2688 6264 2752
rect 6328 2688 6344 2752
rect 6408 2688 6424 2752
rect 6488 2688 6496 2752
rect 6176 2128 6496 2688
rect 6836 8186 7156 8228
rect 6836 7950 6878 8186
rect 7114 7950 7156 8186
rect 6836 7648 7156 7950
rect 6836 7584 6844 7648
rect 6908 7584 6924 7648
rect 6988 7584 7004 7648
rect 7068 7584 7084 7648
rect 7148 7584 7156 7648
rect 6836 6691 7156 7584
rect 6836 6560 6878 6691
rect 7114 6560 7156 6691
rect 6836 6496 6844 6560
rect 7148 6496 7156 6560
rect 6836 6455 6878 6496
rect 7114 6455 7156 6496
rect 6836 5472 7156 6455
rect 6836 5408 6844 5472
rect 6908 5408 6924 5472
rect 6988 5408 7004 5472
rect 7068 5408 7084 5472
rect 7148 5408 7156 5472
rect 6836 5196 7156 5408
rect 6836 4960 6878 5196
rect 7114 4960 7156 5196
rect 6836 4384 7156 4960
rect 6836 4320 6844 4384
rect 6908 4320 6924 4384
rect 6988 4320 7004 4384
rect 7068 4320 7084 4384
rect 7148 4320 7156 4384
rect 6836 3701 7156 4320
rect 6836 3465 6878 3701
rect 7114 3465 7156 3701
rect 6836 3296 7156 3465
rect 6836 3232 6844 3296
rect 6908 3232 6924 3296
rect 6988 3232 7004 3296
rect 7068 3232 7084 3296
rect 7148 3232 7156 3296
rect 6836 2208 7156 3232
rect 6836 2144 6844 2208
rect 6908 2144 6924 2208
rect 6988 2144 7004 2208
rect 7068 2144 7084 2208
rect 7148 2144 7156 2208
rect 6836 2128 7156 2144
<< via4 >>
rect 1733 7290 1969 7526
rect 1733 6016 1969 6031
rect 1733 5952 1763 6016
rect 1763 5952 1779 6016
rect 1779 5952 1843 6016
rect 1843 5952 1859 6016
rect 1859 5952 1923 6016
rect 1923 5952 1939 6016
rect 1939 5952 1969 6016
rect 1733 5795 1969 5952
rect 1733 4300 1969 4536
rect 1733 2805 1969 3041
rect 2393 7950 2629 8186
rect 2393 6560 2629 6691
rect 2393 6496 2423 6560
rect 2423 6496 2439 6560
rect 2439 6496 2503 6560
rect 2503 6496 2519 6560
rect 2519 6496 2583 6560
rect 2583 6496 2599 6560
rect 2599 6496 2629 6560
rect 2393 6455 2629 6496
rect 2393 4960 2629 5196
rect 2393 3465 2629 3701
rect 3228 7290 3464 7526
rect 3228 6016 3464 6031
rect 3228 5952 3258 6016
rect 3258 5952 3274 6016
rect 3274 5952 3338 6016
rect 3338 5952 3354 6016
rect 3354 5952 3418 6016
rect 3418 5952 3434 6016
rect 3434 5952 3464 6016
rect 3228 5795 3464 5952
rect 3228 4300 3464 4536
rect 3228 2805 3464 3041
rect 3888 7950 4124 8186
rect 3888 6560 4124 6691
rect 3888 6496 3918 6560
rect 3918 6496 3934 6560
rect 3934 6496 3998 6560
rect 3998 6496 4014 6560
rect 4014 6496 4078 6560
rect 4078 6496 4094 6560
rect 4094 6496 4124 6560
rect 3888 6455 4124 6496
rect 3888 4960 4124 5196
rect 3888 3465 4124 3701
rect 4723 7290 4959 7526
rect 4723 6016 4959 6031
rect 4723 5952 4753 6016
rect 4753 5952 4769 6016
rect 4769 5952 4833 6016
rect 4833 5952 4849 6016
rect 4849 5952 4913 6016
rect 4913 5952 4929 6016
rect 4929 5952 4959 6016
rect 4723 5795 4959 5952
rect 4723 4300 4959 4536
rect 4723 2805 4959 3041
rect 5383 7950 5619 8186
rect 5383 6560 5619 6691
rect 5383 6496 5413 6560
rect 5413 6496 5429 6560
rect 5429 6496 5493 6560
rect 5493 6496 5509 6560
rect 5509 6496 5573 6560
rect 5573 6496 5589 6560
rect 5589 6496 5619 6560
rect 5383 6455 5619 6496
rect 5383 4960 5619 5196
rect 5383 3465 5619 3701
rect 6218 7290 6454 7526
rect 6218 6016 6454 6031
rect 6218 5952 6248 6016
rect 6248 5952 6264 6016
rect 6264 5952 6328 6016
rect 6328 5952 6344 6016
rect 6344 5952 6408 6016
rect 6408 5952 6424 6016
rect 6424 5952 6454 6016
rect 6218 5795 6454 5952
rect 6218 4300 6454 4536
rect 6218 2805 6454 3041
rect 6878 7950 7114 8186
rect 6878 6560 7114 6691
rect 6878 6496 6908 6560
rect 6908 6496 6924 6560
rect 6924 6496 6988 6560
rect 6988 6496 7004 6560
rect 7004 6496 7068 6560
rect 7068 6496 7084 6560
rect 7084 6496 7114 6560
rect 6878 6455 7114 6496
rect 6878 4960 7114 5196
rect 6878 3465 7114 3701
<< metal5 >>
rect 1056 8186 7156 8228
rect 1056 7950 2393 8186
rect 2629 7950 3888 8186
rect 4124 7950 5383 8186
rect 5619 7950 6878 8186
rect 7114 7950 7156 8186
rect 1056 7908 7156 7950
rect 1056 7526 7132 7568
rect 1056 7290 1733 7526
rect 1969 7290 3228 7526
rect 3464 7290 4723 7526
rect 4959 7290 6218 7526
rect 6454 7290 7132 7526
rect 1056 7248 7132 7290
rect 1056 6691 7156 6733
rect 1056 6455 2393 6691
rect 2629 6455 3888 6691
rect 4124 6455 5383 6691
rect 5619 6455 6878 6691
rect 7114 6455 7156 6691
rect 1056 6413 7156 6455
rect 1056 6031 7132 6073
rect 1056 5795 1733 6031
rect 1969 5795 3228 6031
rect 3464 5795 4723 6031
rect 4959 5795 6218 6031
rect 6454 5795 7132 6031
rect 1056 5753 7132 5795
rect 1056 5196 7156 5238
rect 1056 4960 2393 5196
rect 2629 4960 3888 5196
rect 4124 4960 5383 5196
rect 5619 4960 6878 5196
rect 7114 4960 7156 5196
rect 1056 4918 7156 4960
rect 1056 4536 7132 4578
rect 1056 4300 1733 4536
rect 1969 4300 3228 4536
rect 3464 4300 4723 4536
rect 4959 4300 6218 4536
rect 6454 4300 7132 4536
rect 1056 4258 7132 4300
rect 1056 3701 7156 3743
rect 1056 3465 2393 3701
rect 2629 3465 3888 3701
rect 4124 3465 5383 3701
rect 5619 3465 6878 3701
rect 7114 3465 7156 3701
rect 1056 3423 7156 3465
rect 1056 3041 7132 3083
rect 1056 2805 1733 3041
rect 1969 2805 3228 3041
rect 3464 2805 4723 3041
rect 4959 2805 6218 3041
rect 6454 2805 7132 3041
rect 1056 2763 7132 2805
use sky130_fd_sc_hd__mux2_1  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5060 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _14_
timestamp 1723858470
transform -1 0 2576 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1723858470
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _16_
timestamp 1723858470
transform 1 0 2760 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1723858470
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _18_
timestamp 1723858470
transform 1 0 5612 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1723858470
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _21_
timestamp 1723858470
transform -1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _22_
timestamp 1723858470
transform -1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _23_
timestamp 1723858470
transform -1 0 6164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4232 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _25_
timestamp 1723858470
transform 1 0 2024 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _26_
timestamp 1723858470
transform 1 0 1656 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _27_
timestamp 1723858470
transform 1 0 4784 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1723858470
transform -1 0 3220 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1723858470
transform 1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1723858470
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_33
timestamp 1723858470
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57
timestamp 1723858470
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_26
timestamp 1723858470
transform 1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_34
timestamp 1723858470
transform 1 0 4232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57
timestamp 1723858470
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 1723858470
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1723858470
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 1723858470
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_41
timestamp 1723858470
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_48
timestamp 1723858470
transform 1 0 5520 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_60
timestamp 1723858470
transform 1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1723858470
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_15
timestamp 1723858470
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_26
timestamp 1723858470
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_32
timestamp 1723858470
transform 1 0 4048 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5152 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_57
timestamp 1723858470
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_61
timestamp 1723858470
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 1723858470
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_13
timestamp 1723858470
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_17
timestamp 1723858470
transform 1 0 2668 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1723858470
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_58
timestamp 1723858470
transform 1 0 6440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1723858470
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_30
timestamp 1723858470
transform 1 0 3864 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_34
timestamp 1723858470
transform 1 0 4232 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1723858470
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_57
timestamp 1723858470
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_61
timestamp 1723858470
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_3
timestamp 1723858470
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_16
timestamp 1723858470
transform 1 0 2576 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_29
timestamp 1723858470
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_37
timestamp 1723858470
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_60
timestamp 1723858470
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1723858470
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1723858470
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1723858470
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_39
timestamp 1723858470
transform 1 0 4692 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_57
timestamp 1723858470
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_61
timestamp 1723858470
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1723858470
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1723858470
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1723858470
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1723858470
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_53
timestamp 1723858470
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1723858470
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1723858470
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1723858470
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1723858470
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1723858470
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1723858470
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_57
timestamp 1723858470
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_61
timestamp 1723858470
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 1723858470
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 1723858470
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 1723858470
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_33
timestamp 1723858470
transform 1 0 4140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_45
timestamp 1723858470
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_49
timestamp 1723858470
transform 1 0 5612 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_57
timestamp 1723858470
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_61
timestamp 1723858470
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1723858470
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1723858470
transform -1 0 5060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1723858470
transform -1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1723858470
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1723858470
transform -1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6256 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output5
timestamp 1723858470
transform -1 0 4232 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output6
timestamp 1723858470
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output7
timestamp 1723858470
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1723858470
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1723858470
transform -1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1723858470
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1723858470
transform -1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1723858470
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1723858470
transform -1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1723858470
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1723858470
transform -1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1723858470
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1723858470
transform -1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1723858470
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1723858470
transform -1 0 7084 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1723858470
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1723858470
transform -1 0 7084 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1723858470
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1723858470
transform -1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1723858470
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1723858470
transform -1 0 7084 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1723858470
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1723858470
transform -1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1723858470
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1723858470
transform -1 0 7084 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1723858470
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1723858470
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1723858470
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1723858470
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1723858470
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1723858470
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1723858470
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1723858470
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1723858470
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1723858470
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1723858470
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1723858470
transform 1 0 6256 0 1 7616
box -38 -48 130 592
<< labels >>
flabel metal2 s 7746 9555 7802 10355 0 FreeSans 224 90 0 0 A
port 0 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 B
port 1 nsew signal tristate
flabel metal3 s 7411 5448 8211 5568 0 FreeSans 480 0 0 0 C
port 2 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 D
port 3 nsew signal tristate
flabel metal4 s 2351 2128 2671 8228 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 3846 2128 4166 8228 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 5341 2128 5661 8228 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 6836 2128 7156 8228 0 FreeSans 1920 90 0 0 VGND
port 4 nsew ground bidirectional
flabel metal5 s 1056 3423 7156 3743 0 FreeSans 2560 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal5 s 1056 4918 7156 5238 0 FreeSans 2560 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal5 s 1056 6413 7156 6733 0 FreeSans 2560 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal5 s 1056 7908 7156 8228 0 FreeSans 2560 0 0 0 VGND
port 4 nsew ground bidirectional
flabel metal4 s 1691 2128 2011 8208 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 3186 2128 3506 8208 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 4681 2128 5001 8208 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal4 s 6176 2128 6496 8208 0 FreeSans 1920 90 0 0 VPWR
port 5 nsew power bidirectional
flabel metal5 s 1056 2763 7132 3083 0 FreeSans 2560 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal5 s 1056 4258 7132 4578 0 FreeSans 2560 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal5 s 1056 5753 7132 6073 0 FreeSans 2560 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal5 s 1056 7248 7132 7568 0 FreeSans 2560 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clk
port 6 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 d_in
port 7 nsew signal input
flabel metal2 s 3238 9555 3294 10355 0 FreeSans 224 90 0 0 en
port 8 nsew signal input
flabel metal3 s 7411 688 8211 808 0 FreeSans 480 0 0 0 rst
port 9 nsew signal input
rlabel via1 4130 7616 4130 7616 0 VGND
rlabel metal1 4094 8160 4094 8160 0 VPWR
rlabel metal1 6900 8058 6900 8058 0 A
rlabel metal2 4554 1095 4554 1095 0 B
rlabel metal1 6716 4046 6716 4046 0 C
rlabel metal3 820 4828 820 4828 0 D
rlabel metal1 5566 3366 5566 3366 0 _00_
rlabel metal1 3818 4250 3818 4250 0 _01_
rlabel metal2 3358 3298 3358 3298 0 _02_
rlabel metal1 6072 5338 6072 5338 0 _03_
rlabel metal2 4554 2856 4554 2856 0 _04_
rlabel metal1 2162 4794 2162 4794 0 _05_
rlabel metal1 1978 3400 1978 3400 0 _06_
rlabel metal1 5329 5882 5329 5882 0 _07_
rlabel metal1 5198 5338 5198 5338 0 _08_
rlabel metal2 2254 5066 2254 5066 0 _09_
rlabel metal1 1794 4624 1794 4624 0 _10_
rlabel metal1 4830 3536 4830 3536 0 _11_
rlabel metal2 46 1843 46 1843 0 clk
rlabel metal1 4784 3094 4784 3094 0 clknet_0_clk
rlabel metal1 1886 3570 1886 3570 0 clknet_1_0__leaf_clk
rlabel metal1 5474 3162 5474 3162 0 clknet_1_1__leaf_clk
rlabel metal3 843 9588 843 9588 0 d_in
rlabel metal1 3772 7854 3772 7854 0 en
rlabel metal1 1840 7718 1840 7718 0 net1
rlabel metal1 5244 4998 5244 4998 0 net10
rlabel metal2 2806 4930 2806 4930 0 net11
rlabel metal1 5750 5134 5750 5134 0 net2
rlabel metal1 5290 3468 5290 3468 0 net3
rlabel metal1 6394 6834 6394 6834 0 net4
rlabel metal2 6026 3536 6026 3536 0 net5
rlabel metal1 4370 5134 4370 5134 0 net6
rlabel metal1 3174 4114 3174 4114 0 net7
rlabel metal1 5290 5202 5290 5202 0 net8
rlabel metal1 6072 6290 6072 6290 0 net9
rlabel metal1 6946 2346 6946 2346 0 rst
<< properties >>
string FIXED_BBOX 0 0 8211 10355
<< end >>
